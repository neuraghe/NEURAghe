VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO U2DKTabstractName STRING ;
END PROPERTYDEFINITIONS

MACRO vbbgen_PULPV3_weakdriver
  CLASS CORE ;
  ORIGIN 0 -0.403 ;
  FOREIGN vbbgen_PULPV3_weakdriver 0 0.403 ;
  SIZE 86.44 BY 40.899 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD1V8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER B1 ;
        RECT 56.708 5.261 71.919 9.732 ;
        RECT 67.419 0.72 71.919 27.79 ;
        RECT 67.419 0.721 86.39 5.221 ;
    END
  END VDD1V8
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER B1 ;
        RECT 0.054 0.721 4.554 25.79 ;
        RECT 0.054 0.721 40.888 5.221 ;
        RECT 36.388 0.72 40.888 13.816 ;
        RECT 34.527 9.316 42.661 13.816 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER B1 ;
        RECT 0.001 29.497 4.501 40.884 ;
        RECT 36.388 14.619 40.888 33.998 ;
        RECT 0.001 29.498 40.889 33.998 ;
        RECT 34.527 14.619 42.661 19.119 ;
    END
  END VDD
  PIN pwell
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER B1 ;
        RECT 44.181 12.259 48.681 40.884 ;
        RECT 6.476 36.384 48.681 40.884 ;
        RECT 44.181 12.259 50.949 16.196 ;
    END
  END pwell
  PIN selP1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.218 0.403 57.278 0.806 ;
    END
  END selP1
  PIN selP0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.018 0.403 57.078 0.806 ;
    END
  END selP0
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.418 0.403 57.478 0.806 ;
    END
  END clk
  PIN selN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 56.618 0.403 56.678 0.806 ;
    END
  END selN0
  PIN selN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 56.818 0.403 56.878 0.806 ;
    END
  END selN1
  PIN nwell
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER B1 ;
        RECT 51.587 6.207 56.087 19.211 ;
        RECT 53.975 12.254 58.475 40.884 ;
        RECT 53.975 36.384 86.386 40.884 ;
    END
  END nwell
  OBS
    LAYER M1 ;
      RECT 0.087 20.696 0.821 40.63 ;
      RECT 0.087 8.41 0.821 18.344 ;
      RECT 0.087 8.41 0.269 20.352 ;
      RECT 0.373 7.758 1.337 7.927 ;
      RECT 1.098 29.586 27.396 40.867 ;
      RECT 1.422 0.72 27.396 41.094 ;
      RECT 27.674 30.902 27.724 40.884 ;
      RECT 27.674 0.811 27.724 20.793 ;
      RECT 27.964 0.811 28.014 20.793 ;
      RECT 27.964 30.902 28.764 40.884 ;
      RECT 28.978 20.903 29.231 40.885 ;
      RECT 29.471 20.903 29.521 40.885 ;
      RECT 29.711 40.642 29.761 41.141 ;
      RECT 27.574 41.091 29.761 41.141 ;
      RECT 27.574 41.075 28.524 41.157 ;
      RECT 29.847 20.72 43.021 41.094 ;
      RECT 28.932 0.72 53.306 11.974 ;
      RECT 53.579 0.834 56.424 0.943 ;
      RECT 53.579 0.834 54.926 0.968 ;
      RECT 53.579 0.834 53.916 5.346 ;
      RECT 43.419 20.72 56.593 41.094 ;
      RECT 56.919 20.903 56.969 40.885 ;
      RECT 57.209 20.903 57.462 40.885 ;
      RECT 57.676 30.902 58.476 40.884 ;
      RECT 58.426 0.811 58.476 20.793 ;
      RECT 58.716 30.902 58.766 40.884 ;
      RECT 58.716 0.811 58.766 20.793 ;
      RECT 56.679 40.642 56.729 41.141 ;
      RECT 56.679 41.091 58.866 41.141 ;
      RECT 57.916 41.075 58.866 41.157 ;
      RECT 59.044 29.586 85.342 40.867 ;
      RECT 59.044 0.72 85.018 41.094 ;
      RECT 85.103 7.758 86.067 7.927 ;
      RECT 85.619 20.696 86.353 40.63 ;
      RECT 85.619 8.41 86.353 18.344 ;
      RECT 86.171 8.41 86.353 20.352 ;
    LAYER M1 SPACING 0.05 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER V1 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER M2 ;
      RECT 0.087 20.696 0.821 40.63 ;
      RECT 0.087 8.41 0.821 18.344 ;
      RECT 1.094 40.787 27.396 40.867 ;
      RECT 1.422 0.72 27.396 41.094 ;
      RECT 27.997 30.926 28.731 40.86 ;
      RECT 28.909 30.387 29.019 41.094 ;
      RECT 29.847 20.72 43.021 41.094 ;
      RECT 28.909 40.984 43.021 41.094 ;
      RECT 28.932 0.72 53.306 11.974 ;
      RECT 53.579 0.834 53.916 5.346 ;
      RECT 56.818 0.403 56.878 13.833 ;
      RECT 57.018 0.403 57.078 15.237 ;
      RECT 57.218 0.403 57.278 15.685 ;
      RECT 57.418 0.403 57.478 16.437 ;
      RECT 43.419 20.72 56.593 41.094 ;
      RECT 57.421 30.387 57.531 41.094 ;
      RECT 43.419 40.984 57.531 41.094 ;
      RECT 57.709 30.926 58.443 40.86 ;
      RECT 59.044 40.787 85.346 40.867 ;
      RECT 59.044 0.72 85.018 41.094 ;
      RECT 85.619 20.696 86.353 40.63 ;
      RECT 85.619 8.41 86.353 18.344 ;
    LAYER M2 SPACING 0.05 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER V2 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER M3 ;
      RECT 0.087 20.696 0.821 40.63 ;
      RECT 0.087 8.41 0.821 18.344 ;
      RECT 1.422 0.72 27.396 41.094 ;
      RECT 27.997 30.926 28.731 40.86 ;
      RECT 29.847 20.72 43.021 41.094 ;
      RECT 28.932 0.72 53.306 11.974 ;
      RECT 43.419 20.72 56.593 41.094 ;
      RECT 56.823 0.423 56.873 0.787 ;
      RECT 57.023 0.423 57.073 0.787 ;
      RECT 57.223 0.423 57.273 0.787 ;
      RECT 57.423 0.423 57.473 0.787 ;
      RECT 57.709 30.926 58.443 40.86 ;
      RECT 59.044 0.72 85.018 41.094 ;
      RECT 85.619 20.696 86.353 40.63 ;
      RECT 85.619 8.41 86.353 18.344 ;
    LAYER M3 SPACING 0.05 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER V3 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER M4 ;
      RECT 0.087 20.696 0.821 40.63 ;
      RECT 0.087 8.41 0.821 18.344 ;
      RECT 1.422 0.72 27.396 41.094 ;
      RECT 27.997 30.926 28.731 40.86 ;
      RECT 29.847 20.72 43.021 41.094 ;
      RECT 28.932 0.72 53.306 11.974 ;
      RECT 53.579 0.834 53.916 13.833 ;
      RECT 54.485 0.834 56.526 0.894 ;
      RECT 54.485 0.834 54.545 1.185 ;
      RECT 43.419 20.72 56.593 41.094 ;
      RECT 57.709 30.926 58.443 40.86 ;
      RECT 57.709 0.909 58.443 20.843 ;
      RECT 59.044 0.72 85.018 41.094 ;
      RECT 85.619 20.696 86.353 40.63 ;
      RECT 85.619 8.41 86.353 18.344 ;
    LAYER M4 SPACING 0.05 ;
      RECT 0 0.403 56.526 41.302 ;
      RECT 57.57 0.403 86.44 41.302 ;
      RECT 0 0.898 86.44 41.302 ;
    LAYER M5 ;
      RECT 0.087 20.696 0.821 40.63 ;
      RECT 0.087 8.41 0.821 18.344 ;
      RECT 1.422 0.72 27.396 41.094 ;
      RECT 27.997 30.926 28.731 40.86 ;
      RECT 29.847 20.72 43.021 41.094 ;
      RECT 28.932 0.72 53.306 11.974 ;
      RECT 43.419 20.72 56.593 41.094 ;
      RECT 57.709 30.926 58.443 40.86 ;
      RECT 57.709 0.909 58.443 20.843 ;
      RECT 59.044 0.72 85.018 41.094 ;
      RECT 85.619 20.696 86.353 40.63 ;
      RECT 85.619 8.41 86.353 18.344 ;
    LAYER M5 SPACING 0.05 ;
      RECT 0 0.403 56.511 41.302 ;
      RECT 57.585 0.403 86.44 41.302 ;
      RECT 0 0.913 86.44 41.302 ;
    LAYER M6 ;
      RECT 0.054 8.386 2.554 18.368 ;
      RECT 0.054 23.29 18.939 25.79 ;
      RECT 0.054 29.249 17.151 31.749 ;
      RECT 0.054 35.272 16.586 37.772 ;
      RECT 0.054 20.671 2.554 40.654 ;
      RECT 27.964 30.902 30.464 40.884 ;
      RECT 55.976 30.902 58.476 40.884 ;
      RECT 27.964 36.384 58.476 40.884 ;
      RECT 14.521 0.72 71.919 3.22 ;
      RECT 14.521 0.72 19.021 18.368 ;
      RECT 67.419 0.72 71.919 18.368 ;
      RECT 67.501 23.29 86.386 25.79 ;
      RECT 69.289 29.249 86.386 31.749 ;
      RECT 69.854 35.272 86.386 37.772 ;
      RECT 83.886 20.671 86.386 40.654 ;
      RECT 83.886 8.386 86.386 18.368 ;
    LAYER M6 SPACING 0.05 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER V4 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER V5 ;
      RECT 0 0.403 86.44 41.302 ;
    LAYER W0 ;
      RECT 17.986 3.075 18.086 3.175 ;
      RECT 17.986 2.745 18.086 2.845 ;
      RECT 17.986 2.415 18.086 2.515 ;
      RECT 17.986 2.085 18.086 2.185 ;
      RECT 17.986 1.755 18.086 1.855 ;
      RECT 17.986 1.425 18.086 1.525 ;
      RECT 17.986 1.095 18.086 1.195 ;
      RECT 17.986 0.765 18.086 0.865 ;
      RECT 18.316 3.075 18.416 3.175 ;
      RECT 18.316 2.745 18.416 2.845 ;
      RECT 18.316 2.415 18.416 2.515 ;
      RECT 18.316 2.085 18.416 2.185 ;
      RECT 18.316 1.755 18.416 1.855 ;
      RECT 18.316 1.425 18.416 1.525 ;
      RECT 18.316 1.095 18.416 1.195 ;
      RECT 18.316 0.765 18.416 0.865 ;
      RECT 18.646 3.075 18.746 3.175 ;
      RECT 18.646 2.745 18.746 2.845 ;
      RECT 18.646 2.415 18.746 2.515 ;
      RECT 18.646 2.085 18.746 2.185 ;
      RECT 18.646 1.755 18.746 1.855 ;
      RECT 18.646 1.425 18.746 1.525 ;
      RECT 18.646 1.095 18.746 1.195 ;
      RECT 18.646 0.765 18.746 0.865 ;
      RECT 18.976 3.075 19.076 3.175 ;
      RECT 18.976 2.745 19.076 2.845 ;
      RECT 18.976 2.415 19.076 2.515 ;
      RECT 18.976 2.085 19.076 2.185 ;
      RECT 18.976 1.755 19.076 1.855 ;
      RECT 18.976 1.425 19.076 1.525 ;
      RECT 18.976 1.095 19.076 1.195 ;
      RECT 18.976 0.765 19.076 0.865 ;
      RECT 19.306 3.075 19.406 3.175 ;
      RECT 19.306 2.745 19.406 2.845 ;
      RECT 19.306 2.415 19.406 2.515 ;
      RECT 19.306 2.085 19.406 2.185 ;
      RECT 19.306 1.755 19.406 1.855 ;
      RECT 19.306 1.425 19.406 1.525 ;
      RECT 19.306 1.095 19.406 1.195 ;
      RECT 19.306 0.765 19.406 0.865 ;
      RECT 19.636 3.075 19.736 3.175 ;
      RECT 19.636 2.745 19.736 2.845 ;
      RECT 19.636 2.415 19.736 2.515 ;
      RECT 19.636 2.085 19.736 2.185 ;
      RECT 19.636 1.755 19.736 1.855 ;
      RECT 19.636 1.425 19.736 1.525 ;
      RECT 19.636 1.095 19.736 1.195 ;
      RECT 19.636 0.765 19.736 0.865 ;
      RECT 19.966 3.075 20.066 3.175 ;
      RECT 19.966 2.745 20.066 2.845 ;
      RECT 19.966 2.415 20.066 2.515 ;
      RECT 19.966 2.085 20.066 2.185 ;
      RECT 19.966 1.755 20.066 1.855 ;
      RECT 19.966 1.425 20.066 1.525 ;
      RECT 19.966 1.095 20.066 1.195 ;
      RECT 19.966 0.765 20.066 0.865 ;
      RECT 20.296 3.075 20.396 3.175 ;
      RECT 20.296 2.745 20.396 2.845 ;
      RECT 20.296 2.415 20.396 2.515 ;
      RECT 20.296 2.085 20.396 2.185 ;
      RECT 20.296 1.755 20.396 1.855 ;
      RECT 20.296 1.425 20.396 1.525 ;
      RECT 20.296 1.095 20.396 1.195 ;
      RECT 20.296 0.765 20.396 0.865 ;
      RECT 20.626 3.075 20.726 3.175 ;
      RECT 20.626 2.745 20.726 2.845 ;
      RECT 20.626 2.415 20.726 2.515 ;
      RECT 20.626 2.085 20.726 2.185 ;
      RECT 20.626 1.755 20.726 1.855 ;
      RECT 20.626 1.425 20.726 1.525 ;
      RECT 20.626 1.095 20.726 1.195 ;
      RECT 20.626 0.765 20.726 0.865 ;
      RECT 20.956 3.075 21.056 3.175 ;
      RECT 20.956 2.745 21.056 2.845 ;
      RECT 20.956 2.415 21.056 2.515 ;
      RECT 20.956 2.085 21.056 2.185 ;
      RECT 20.956 1.755 21.056 1.855 ;
      RECT 20.956 1.425 21.056 1.525 ;
      RECT 20.956 1.095 21.056 1.195 ;
      RECT 20.956 0.765 21.056 0.865 ;
      RECT 21.286 3.075 21.386 3.175 ;
      RECT 21.286 2.745 21.386 2.845 ;
      RECT 21.286 2.415 21.386 2.515 ;
      RECT 21.286 2.085 21.386 2.185 ;
      RECT 21.286 1.755 21.386 1.855 ;
      RECT 21.286 1.425 21.386 1.525 ;
      RECT 21.286 1.095 21.386 1.195 ;
      RECT 21.286 0.765 21.386 0.865 ;
      RECT 21.616 3.075 21.716 3.175 ;
      RECT 21.616 2.745 21.716 2.845 ;
      RECT 21.616 2.415 21.716 2.515 ;
      RECT 21.616 2.085 21.716 2.185 ;
      RECT 21.616 1.755 21.716 1.855 ;
      RECT 21.616 1.425 21.716 1.525 ;
      RECT 21.616 1.095 21.716 1.195 ;
      RECT 21.616 0.765 21.716 0.865 ;
      RECT 21.946 3.075 22.046 3.175 ;
      RECT 21.946 2.745 22.046 2.845 ;
      RECT 21.946 2.415 22.046 2.515 ;
      RECT 21.946 2.085 22.046 2.185 ;
      RECT 21.946 1.755 22.046 1.855 ;
      RECT 21.946 1.425 22.046 1.525 ;
      RECT 21.946 1.095 22.046 1.195 ;
      RECT 21.946 0.765 22.046 0.865 ;
      RECT 22.276 3.075 22.376 3.175 ;
      RECT 22.276 2.745 22.376 2.845 ;
      RECT 22.276 2.415 22.376 2.515 ;
      RECT 22.276 2.085 22.376 2.185 ;
      RECT 22.276 1.755 22.376 1.855 ;
      RECT 22.276 1.425 22.376 1.525 ;
      RECT 22.276 1.095 22.376 1.195 ;
      RECT 22.276 0.765 22.376 0.865 ;
      RECT 22.606 3.075 22.706 3.175 ;
      RECT 22.606 2.745 22.706 2.845 ;
      RECT 22.606 2.415 22.706 2.515 ;
      RECT 22.606 2.085 22.706 2.185 ;
      RECT 22.606 1.755 22.706 1.855 ;
      RECT 22.606 1.425 22.706 1.525 ;
      RECT 22.606 1.095 22.706 1.195 ;
      RECT 22.606 0.765 22.706 0.865 ;
      RECT 22.936 3.075 23.036 3.175 ;
      RECT 22.936 2.745 23.036 2.845 ;
      RECT 22.936 2.415 23.036 2.515 ;
      RECT 22.936 2.085 23.036 2.185 ;
      RECT 22.936 1.755 23.036 1.855 ;
      RECT 22.936 1.425 23.036 1.525 ;
      RECT 22.936 1.095 23.036 1.195 ;
      RECT 22.936 0.765 23.036 0.865 ;
      RECT 23.266 3.075 23.366 3.175 ;
      RECT 23.266 2.745 23.366 2.845 ;
      RECT 23.266 2.415 23.366 2.515 ;
      RECT 23.266 2.085 23.366 2.185 ;
      RECT 23.266 1.755 23.366 1.855 ;
      RECT 23.266 1.425 23.366 1.525 ;
      RECT 23.266 1.095 23.366 1.195 ;
      RECT 23.266 0.765 23.366 0.865 ;
      RECT 23.596 3.075 23.696 3.175 ;
      RECT 23.596 2.745 23.696 2.845 ;
      RECT 23.596 2.415 23.696 2.515 ;
      RECT 23.596 2.085 23.696 2.185 ;
      RECT 23.596 1.755 23.696 1.855 ;
      RECT 23.596 1.425 23.696 1.525 ;
      RECT 23.596 1.095 23.696 1.195 ;
      RECT 23.596 0.765 23.696 0.865 ;
      RECT 23.926 3.075 24.026 3.175 ;
      RECT 23.926 2.745 24.026 2.845 ;
      RECT 23.926 2.415 24.026 2.515 ;
      RECT 23.926 2.085 24.026 2.185 ;
      RECT 23.926 1.755 24.026 1.855 ;
      RECT 23.926 1.425 24.026 1.525 ;
      RECT 23.926 1.095 24.026 1.195 ;
      RECT 23.926 0.765 24.026 0.865 ;
      RECT 24.256 3.075 24.356 3.175 ;
      RECT 24.256 2.745 24.356 2.845 ;
      RECT 24.256 2.415 24.356 2.515 ;
      RECT 24.256 2.085 24.356 2.185 ;
      RECT 24.256 1.755 24.356 1.855 ;
      RECT 24.256 1.425 24.356 1.525 ;
      RECT 24.256 1.095 24.356 1.195 ;
      RECT 24.256 0.765 24.356 0.865 ;
      RECT 24.586 3.075 24.686 3.175 ;
      RECT 24.586 2.745 24.686 2.845 ;
      RECT 24.586 2.415 24.686 2.515 ;
      RECT 24.586 2.085 24.686 2.185 ;
      RECT 24.586 1.755 24.686 1.855 ;
      RECT 24.586 1.425 24.686 1.525 ;
      RECT 24.586 1.095 24.686 1.195 ;
      RECT 24.586 0.765 24.686 0.865 ;
      RECT 24.916 3.075 25.016 3.175 ;
      RECT 24.916 2.745 25.016 2.845 ;
      RECT 24.916 2.415 25.016 2.515 ;
      RECT 24.916 2.085 25.016 2.185 ;
      RECT 24.916 1.755 25.016 1.855 ;
      RECT 24.916 1.425 25.016 1.525 ;
      RECT 24.916 1.095 25.016 1.195 ;
      RECT 24.916 0.765 25.016 0.865 ;
      RECT 25.246 3.075 25.346 3.175 ;
      RECT 25.246 2.745 25.346 2.845 ;
      RECT 25.246 2.415 25.346 2.515 ;
      RECT 25.246 2.085 25.346 2.185 ;
      RECT 25.246 1.755 25.346 1.855 ;
      RECT 25.246 1.425 25.346 1.525 ;
      RECT 25.246 1.095 25.346 1.195 ;
      RECT 25.246 0.765 25.346 0.865 ;
      RECT 25.576 3.075 25.676 3.175 ;
      RECT 25.576 2.745 25.676 2.845 ;
      RECT 25.576 2.415 25.676 2.515 ;
      RECT 25.576 2.085 25.676 2.185 ;
      RECT 25.576 1.755 25.676 1.855 ;
      RECT 25.576 1.425 25.676 1.525 ;
      RECT 25.576 1.095 25.676 1.195 ;
      RECT 25.576 0.765 25.676 0.865 ;
      RECT 25.906 3.075 26.006 3.175 ;
      RECT 25.906 2.745 26.006 2.845 ;
      RECT 25.906 2.415 26.006 2.515 ;
      RECT 25.906 2.085 26.006 2.185 ;
      RECT 25.906 1.755 26.006 1.855 ;
      RECT 25.906 1.425 26.006 1.525 ;
      RECT 25.906 1.095 26.006 1.195 ;
      RECT 25.906 0.765 26.006 0.865 ;
      RECT 26.236 3.075 26.336 3.175 ;
      RECT 26.236 2.745 26.336 2.845 ;
      RECT 26.236 2.415 26.336 2.515 ;
      RECT 26.236 2.085 26.336 2.185 ;
      RECT 26.236 1.755 26.336 1.855 ;
      RECT 26.236 1.425 26.336 1.525 ;
      RECT 26.236 1.095 26.336 1.195 ;
      RECT 26.236 0.765 26.336 0.865 ;
      RECT 26.566 3.075 26.666 3.175 ;
      RECT 26.566 2.745 26.666 2.845 ;
      RECT 26.566 2.415 26.666 2.515 ;
      RECT 26.566 2.085 26.666 2.185 ;
      RECT 26.566 1.755 26.666 1.855 ;
      RECT 26.566 1.425 26.666 1.525 ;
      RECT 26.566 1.095 26.666 1.195 ;
      RECT 26.566 0.765 26.666 0.865 ;
      RECT 26.896 3.075 26.996 3.175 ;
      RECT 26.896 2.745 26.996 2.845 ;
      RECT 26.896 2.415 26.996 2.515 ;
      RECT 26.896 2.085 26.996 2.185 ;
      RECT 26.896 1.755 26.996 1.855 ;
      RECT 26.896 1.425 26.996 1.525 ;
      RECT 26.896 1.095 26.996 1.195 ;
      RECT 26.896 0.765 26.996 0.865 ;
      RECT 27.226 3.075 27.326 3.175 ;
      RECT 27.226 2.745 27.326 2.845 ;
      RECT 27.226 2.415 27.326 2.515 ;
      RECT 27.226 2.085 27.326 2.185 ;
      RECT 27.226 1.755 27.326 1.855 ;
      RECT 27.226 1.425 27.326 1.525 ;
      RECT 27.226 1.095 27.326 1.195 ;
      RECT 27.226 0.765 27.326 0.865 ;
      RECT 27.556 3.075 27.656 3.175 ;
      RECT 27.556 2.745 27.656 2.845 ;
      RECT 27.556 2.415 27.656 2.515 ;
      RECT 27.556 2.085 27.656 2.185 ;
      RECT 27.556 1.755 27.656 1.855 ;
      RECT 27.556 1.425 27.656 1.525 ;
      RECT 27.556 1.095 27.656 1.195 ;
      RECT 27.556 0.765 27.656 0.865 ;
      RECT 27.886 3.075 27.986 3.175 ;
      RECT 27.886 2.745 27.986 2.845 ;
      RECT 27.886 2.415 27.986 2.515 ;
      RECT 27.886 2.085 27.986 2.185 ;
      RECT 27.886 1.755 27.986 1.855 ;
      RECT 27.886 1.425 27.986 1.525 ;
      RECT 27.886 1.095 27.986 1.195 ;
      RECT 27.886 0.765 27.986 0.865 ;
      RECT 28.216 3.075 28.316 3.175 ;
      RECT 28.216 2.745 28.316 2.845 ;
      RECT 28.216 2.415 28.316 2.515 ;
      RECT 28.216 2.085 28.316 2.185 ;
      RECT 28.216 1.755 28.316 1.855 ;
      RECT 28.216 1.425 28.316 1.525 ;
      RECT 28.216 1.095 28.316 1.195 ;
      RECT 28.216 0.765 28.316 0.865 ;
      RECT 28.546 3.075 28.646 3.175 ;
      RECT 28.546 2.745 28.646 2.845 ;
      RECT 28.546 2.415 28.646 2.515 ;
      RECT 28.546 2.085 28.646 2.185 ;
      RECT 28.546 1.755 28.646 1.855 ;
      RECT 28.546 1.425 28.646 1.525 ;
      RECT 28.546 1.095 28.646 1.195 ;
      RECT 28.546 0.765 28.646 0.865 ;
      RECT 28.876 3.075 28.976 3.175 ;
      RECT 28.876 2.745 28.976 2.845 ;
      RECT 28.876 2.415 28.976 2.515 ;
      RECT 28.876 2.085 28.976 2.185 ;
      RECT 28.876 1.755 28.976 1.855 ;
      RECT 28.876 1.425 28.976 1.525 ;
      RECT 28.876 1.095 28.976 1.195 ;
      RECT 28.876 0.765 28.976 0.865 ;
      RECT 29.206 3.075 29.306 3.175 ;
      RECT 29.206 2.745 29.306 2.845 ;
      RECT 29.206 2.415 29.306 2.515 ;
      RECT 29.206 2.085 29.306 2.185 ;
      RECT 29.206 1.755 29.306 1.855 ;
      RECT 29.206 1.425 29.306 1.525 ;
      RECT 29.206 1.095 29.306 1.195 ;
      RECT 29.206 0.765 29.306 0.865 ;
      RECT 29.536 3.075 29.636 3.175 ;
      RECT 29.536 2.745 29.636 2.845 ;
      RECT 29.536 2.415 29.636 2.515 ;
      RECT 29.536 2.085 29.636 2.185 ;
      RECT 29.536 1.755 29.636 1.855 ;
      RECT 29.536 1.425 29.636 1.525 ;
      RECT 29.536 1.095 29.636 1.195 ;
      RECT 29.536 0.765 29.636 0.865 ;
      RECT 29.866 3.075 29.966 3.175 ;
      RECT 29.866 2.745 29.966 2.845 ;
      RECT 29.866 2.415 29.966 2.515 ;
      RECT 29.866 2.085 29.966 2.185 ;
      RECT 29.866 1.755 29.966 1.855 ;
      RECT 29.866 1.425 29.966 1.525 ;
      RECT 29.866 1.095 29.966 1.195 ;
      RECT 29.866 0.765 29.966 0.865 ;
      RECT 30.196 3.075 30.296 3.175 ;
      RECT 30.196 2.745 30.296 2.845 ;
      RECT 30.196 2.415 30.296 2.515 ;
      RECT 30.196 2.085 30.296 2.185 ;
      RECT 30.196 1.755 30.296 1.855 ;
      RECT 30.196 1.425 30.296 1.525 ;
      RECT 30.196 1.095 30.296 1.195 ;
      RECT 30.196 0.765 30.296 0.865 ;
      RECT 30.526 3.075 30.626 3.175 ;
      RECT 30.526 2.745 30.626 2.845 ;
      RECT 30.526 2.415 30.626 2.515 ;
      RECT 30.526 2.085 30.626 2.185 ;
      RECT 30.526 1.755 30.626 1.855 ;
      RECT 30.526 1.425 30.626 1.525 ;
      RECT 30.526 1.095 30.626 1.195 ;
      RECT 30.526 0.765 30.626 0.865 ;
      RECT 30.856 3.075 30.956 3.175 ;
      RECT 30.856 2.745 30.956 2.845 ;
      RECT 30.856 2.415 30.956 2.515 ;
      RECT 30.856 2.085 30.956 2.185 ;
      RECT 30.856 1.755 30.956 1.855 ;
      RECT 30.856 1.425 30.956 1.525 ;
      RECT 30.856 1.095 30.956 1.195 ;
      RECT 30.856 0.765 30.956 0.865 ;
      RECT 31.186 3.075 31.286 3.175 ;
      RECT 31.186 2.745 31.286 2.845 ;
      RECT 31.186 2.415 31.286 2.515 ;
      RECT 31.186 2.085 31.286 2.185 ;
      RECT 31.186 1.755 31.286 1.855 ;
      RECT 31.186 1.425 31.286 1.525 ;
      RECT 31.186 1.095 31.286 1.195 ;
      RECT 31.186 0.765 31.286 0.865 ;
      RECT 31.516 3.075 31.616 3.175 ;
      RECT 31.516 2.745 31.616 2.845 ;
      RECT 31.516 2.415 31.616 2.515 ;
      RECT 31.516 2.085 31.616 2.185 ;
      RECT 31.516 1.755 31.616 1.855 ;
      RECT 31.516 1.425 31.616 1.525 ;
      RECT 31.516 1.095 31.616 1.195 ;
      RECT 31.516 0.765 31.616 0.865 ;
      RECT 31.846 3.075 31.946 3.175 ;
      RECT 31.846 2.745 31.946 2.845 ;
      RECT 31.846 2.415 31.946 2.515 ;
      RECT 31.846 2.085 31.946 2.185 ;
      RECT 31.846 1.755 31.946 1.855 ;
      RECT 31.846 1.425 31.946 1.525 ;
      RECT 31.846 1.095 31.946 1.195 ;
      RECT 31.846 0.765 31.946 0.865 ;
      RECT 32.176 3.075 32.276 3.175 ;
      RECT 32.176 2.745 32.276 2.845 ;
      RECT 32.176 2.415 32.276 2.515 ;
      RECT 32.176 2.085 32.276 2.185 ;
      RECT 32.176 1.755 32.276 1.855 ;
      RECT 32.176 1.425 32.276 1.525 ;
      RECT 32.176 1.095 32.276 1.195 ;
      RECT 32.176 0.765 32.276 0.865 ;
      RECT 32.324 25.968 32.424 26.068 ;
      RECT 32.324 25.638 32.424 25.738 ;
      RECT 32.324 25.308 32.424 25.408 ;
      RECT 32.324 24.978 32.424 25.078 ;
      RECT 32.324 24.648 32.424 24.748 ;
      RECT 32.324 24.318 32.424 24.418 ;
      RECT 32.324 23.988 32.424 24.088 ;
      RECT 32.324 23.658 32.424 23.758 ;
      RECT 32.324 23.328 32.424 23.428 ;
      RECT 32.324 13.35 32.424 13.45 ;
      RECT 32.324 13.02 32.424 13.12 ;
      RECT 32.506 3.075 32.606 3.175 ;
      RECT 32.506 2.745 32.606 2.845 ;
      RECT 32.506 2.415 32.606 2.515 ;
      RECT 32.506 2.085 32.606 2.185 ;
      RECT 32.506 1.755 32.606 1.855 ;
      RECT 32.506 1.425 32.606 1.525 ;
      RECT 32.506 1.095 32.606 1.195 ;
      RECT 32.506 0.765 32.606 0.865 ;
      RECT 32.654 25.968 32.754 26.068 ;
      RECT 32.654 25.638 32.754 25.738 ;
      RECT 32.654 25.308 32.754 25.408 ;
      RECT 32.654 24.978 32.754 25.078 ;
      RECT 32.654 24.648 32.754 24.748 ;
      RECT 32.654 24.318 32.754 24.418 ;
      RECT 32.654 23.988 32.754 24.088 ;
      RECT 32.654 23.658 32.754 23.758 ;
      RECT 32.654 23.328 32.754 23.428 ;
      RECT 32.654 13.35 32.754 13.45 ;
      RECT 32.654 13.02 32.754 13.12 ;
      RECT 32.836 3.075 32.936 3.175 ;
      RECT 32.836 2.745 32.936 2.845 ;
      RECT 32.836 2.415 32.936 2.515 ;
      RECT 32.836 2.085 32.936 2.185 ;
      RECT 32.836 1.755 32.936 1.855 ;
      RECT 32.836 1.425 32.936 1.525 ;
      RECT 32.836 1.095 32.936 1.195 ;
      RECT 32.836 0.765 32.936 0.865 ;
      RECT 32.984 25.968 33.084 26.068 ;
      RECT 32.984 25.638 33.084 25.738 ;
      RECT 32.984 25.308 33.084 25.408 ;
      RECT 32.984 24.978 33.084 25.078 ;
      RECT 32.984 24.648 33.084 24.748 ;
      RECT 32.984 24.318 33.084 24.418 ;
      RECT 32.984 23.988 33.084 24.088 ;
      RECT 32.984 23.658 33.084 23.758 ;
      RECT 32.984 23.328 33.084 23.428 ;
      RECT 32.984 13.35 33.084 13.45 ;
      RECT 32.984 13.02 33.084 13.12 ;
      RECT 33.166 3.075 33.266 3.175 ;
      RECT 33.166 2.745 33.266 2.845 ;
      RECT 33.166 2.415 33.266 2.515 ;
      RECT 33.166 2.085 33.266 2.185 ;
      RECT 33.166 1.755 33.266 1.855 ;
      RECT 33.166 1.425 33.266 1.525 ;
      RECT 33.166 1.095 33.266 1.195 ;
      RECT 33.166 0.765 33.266 0.865 ;
      RECT 33.496 3.075 33.596 3.175 ;
      RECT 33.496 2.745 33.596 2.845 ;
      RECT 33.496 2.415 33.596 2.515 ;
      RECT 33.496 2.085 33.596 2.185 ;
      RECT 33.496 1.755 33.596 1.855 ;
      RECT 33.496 1.425 33.596 1.525 ;
      RECT 33.496 1.095 33.596 1.195 ;
      RECT 33.496 0.765 33.596 0.865 ;
      RECT 33.826 3.075 33.926 3.175 ;
      RECT 33.826 2.745 33.926 2.845 ;
      RECT 33.826 2.415 33.926 2.515 ;
      RECT 33.826 2.085 33.926 2.185 ;
      RECT 33.826 1.755 33.926 1.855 ;
      RECT 33.826 1.425 33.926 1.525 ;
      RECT 33.826 1.095 33.926 1.195 ;
      RECT 33.826 0.765 33.926 0.865 ;
      RECT 34.156 3.075 34.256 3.175 ;
      RECT 34.156 2.745 34.256 2.845 ;
      RECT 34.156 2.415 34.256 2.515 ;
      RECT 34.156 2.085 34.256 2.185 ;
      RECT 34.156 1.755 34.256 1.855 ;
      RECT 34.156 1.425 34.256 1.525 ;
      RECT 34.156 1.095 34.256 1.195 ;
      RECT 34.156 0.765 34.256 0.865 ;
      RECT 34.583 15.51 34.683 15.61 ;
      RECT 34.583 15.18 34.683 15.28 ;
      RECT 34.583 13.12 34.683 13.22 ;
      RECT 34.583 12.79 34.683 12.89 ;
      RECT 34.913 15.51 35.013 15.61 ;
      RECT 34.913 15.18 35.013 15.28 ;
      RECT 34.913 13.12 35.013 13.22 ;
      RECT 34.913 12.79 35.013 12.89 ;
      RECT 35.243 15.51 35.343 15.61 ;
      RECT 35.243 15.18 35.343 15.28 ;
      RECT 35.243 13.12 35.343 13.22 ;
      RECT 35.243 12.79 35.343 12.89 ;
      RECT 35.322 40.729 35.422 40.829 ;
      RECT 35.322 40.399 35.422 40.499 ;
      RECT 35.322 40.069 35.422 40.169 ;
      RECT 35.322 39.739 35.422 39.839 ;
      RECT 35.322 39.409 35.422 39.509 ;
      RECT 35.322 39.079 35.422 39.179 ;
      RECT 35.322 38.749 35.422 38.849 ;
      RECT 35.322 38.419 35.422 38.519 ;
      RECT 35.322 38.089 35.422 38.189 ;
      RECT 35.322 37.759 35.422 37.859 ;
      RECT 35.322 37.429 35.422 37.529 ;
      RECT 35.322 37.099 35.422 37.199 ;
      RECT 35.322 36.769 35.422 36.869 ;
      RECT 35.322 36.439 35.422 36.539 ;
      RECT 35.573 15.51 35.673 15.61 ;
      RECT 35.573 15.18 35.673 15.28 ;
      RECT 35.573 13.12 35.673 13.22 ;
      RECT 35.573 12.79 35.673 12.89 ;
      RECT 35.652 40.729 35.752 40.829 ;
      RECT 35.652 40.399 35.752 40.499 ;
      RECT 35.652 40.069 35.752 40.169 ;
      RECT 35.652 39.739 35.752 39.839 ;
      RECT 35.652 39.409 35.752 39.509 ;
      RECT 35.652 39.079 35.752 39.179 ;
      RECT 35.652 38.749 35.752 38.849 ;
      RECT 35.652 38.419 35.752 38.519 ;
      RECT 35.652 38.089 35.752 38.189 ;
      RECT 35.652 37.759 35.752 37.859 ;
      RECT 35.652 37.429 35.752 37.529 ;
      RECT 35.652 37.099 35.752 37.199 ;
      RECT 35.652 36.769 35.752 36.869 ;
      RECT 35.652 36.439 35.752 36.539 ;
      RECT 35.757 3.075 35.857 3.175 ;
      RECT 35.757 2.745 35.857 2.845 ;
      RECT 35.757 2.415 35.857 2.515 ;
      RECT 35.757 2.085 35.857 2.185 ;
      RECT 35.757 1.755 35.857 1.855 ;
      RECT 35.757 1.425 35.857 1.525 ;
      RECT 35.757 1.095 35.857 1.195 ;
      RECT 35.757 0.765 35.857 0.865 ;
      RECT 35.903 15.51 36.003 15.61 ;
      RECT 35.903 15.18 36.003 15.28 ;
      RECT 35.903 13.12 36.003 13.22 ;
      RECT 35.903 12.79 36.003 12.89 ;
      RECT 35.982 40.729 36.082 40.829 ;
      RECT 35.982 40.399 36.082 40.499 ;
      RECT 35.982 40.069 36.082 40.169 ;
      RECT 35.982 39.739 36.082 39.839 ;
      RECT 35.982 39.409 36.082 39.509 ;
      RECT 35.982 39.079 36.082 39.179 ;
      RECT 35.982 38.749 36.082 38.849 ;
      RECT 35.982 38.419 36.082 38.519 ;
      RECT 35.982 38.089 36.082 38.189 ;
      RECT 35.982 37.759 36.082 37.859 ;
      RECT 35.982 37.429 36.082 37.529 ;
      RECT 35.982 37.099 36.082 37.199 ;
      RECT 35.982 36.769 36.082 36.869 ;
      RECT 35.982 36.439 36.082 36.539 ;
      RECT 36.087 3.075 36.187 3.175 ;
      RECT 36.087 2.745 36.187 2.845 ;
      RECT 36.087 2.415 36.187 2.515 ;
      RECT 36.087 2.085 36.187 2.185 ;
      RECT 36.087 1.755 36.187 1.855 ;
      RECT 36.087 1.425 36.187 1.525 ;
      RECT 36.087 1.095 36.187 1.195 ;
      RECT 36.087 0.765 36.187 0.865 ;
      RECT 36.233 15.51 36.333 15.61 ;
      RECT 36.233 15.18 36.333 15.28 ;
      RECT 36.233 13.12 36.333 13.22 ;
      RECT 36.233 12.79 36.333 12.89 ;
      RECT 36.312 40.729 36.412 40.829 ;
      RECT 36.312 40.399 36.412 40.499 ;
      RECT 36.312 40.069 36.412 40.169 ;
      RECT 36.312 39.739 36.412 39.839 ;
      RECT 36.312 39.409 36.412 39.509 ;
      RECT 36.312 39.079 36.412 39.179 ;
      RECT 36.312 38.749 36.412 38.849 ;
      RECT 36.312 38.419 36.412 38.519 ;
      RECT 36.312 38.089 36.412 38.189 ;
      RECT 36.312 37.759 36.412 37.859 ;
      RECT 36.312 37.429 36.412 37.529 ;
      RECT 36.312 37.099 36.412 37.199 ;
      RECT 36.312 36.769 36.412 36.869 ;
      RECT 36.312 36.439 36.412 36.539 ;
      RECT 36.417 3.075 36.517 3.175 ;
      RECT 36.417 2.745 36.517 2.845 ;
      RECT 36.417 2.415 36.517 2.515 ;
      RECT 36.417 2.085 36.517 2.185 ;
      RECT 36.417 1.755 36.517 1.855 ;
      RECT 36.417 1.425 36.517 1.525 ;
      RECT 36.417 1.095 36.517 1.195 ;
      RECT 36.417 0.765 36.517 0.865 ;
      RECT 36.563 15.51 36.663 15.61 ;
      RECT 36.563 15.18 36.663 15.28 ;
      RECT 36.563 13.12 36.663 13.22 ;
      RECT 36.563 12.79 36.663 12.89 ;
      RECT 36.642 40.729 36.742 40.829 ;
      RECT 36.642 40.399 36.742 40.499 ;
      RECT 36.642 40.069 36.742 40.169 ;
      RECT 36.642 39.739 36.742 39.839 ;
      RECT 36.642 39.409 36.742 39.509 ;
      RECT 36.642 39.079 36.742 39.179 ;
      RECT 36.642 38.749 36.742 38.849 ;
      RECT 36.642 38.419 36.742 38.519 ;
      RECT 36.642 38.089 36.742 38.189 ;
      RECT 36.642 37.759 36.742 37.859 ;
      RECT 36.642 37.429 36.742 37.529 ;
      RECT 36.642 37.099 36.742 37.199 ;
      RECT 36.642 36.769 36.742 36.869 ;
      RECT 36.642 36.439 36.742 36.539 ;
      RECT 36.747 3.075 36.847 3.175 ;
      RECT 36.747 2.745 36.847 2.845 ;
      RECT 36.747 2.415 36.847 2.515 ;
      RECT 36.747 2.085 36.847 2.185 ;
      RECT 36.747 1.755 36.847 1.855 ;
      RECT 36.747 1.425 36.847 1.525 ;
      RECT 36.747 1.095 36.847 1.195 ;
      RECT 36.747 0.765 36.847 0.865 ;
      RECT 36.893 15.51 36.993 15.61 ;
      RECT 36.893 15.18 36.993 15.28 ;
      RECT 36.893 13.12 36.993 13.22 ;
      RECT 36.893 12.79 36.993 12.89 ;
      RECT 36.972 40.729 37.072 40.829 ;
      RECT 36.972 40.399 37.072 40.499 ;
      RECT 36.972 40.069 37.072 40.169 ;
      RECT 36.972 39.739 37.072 39.839 ;
      RECT 36.972 39.409 37.072 39.509 ;
      RECT 36.972 39.079 37.072 39.179 ;
      RECT 36.972 38.749 37.072 38.849 ;
      RECT 36.972 38.419 37.072 38.519 ;
      RECT 36.972 38.089 37.072 38.189 ;
      RECT 36.972 37.759 37.072 37.859 ;
      RECT 36.972 37.429 37.072 37.529 ;
      RECT 36.972 37.099 37.072 37.199 ;
      RECT 36.972 36.769 37.072 36.869 ;
      RECT 36.972 36.439 37.072 36.539 ;
      RECT 37.077 3.075 37.177 3.175 ;
      RECT 37.077 2.745 37.177 2.845 ;
      RECT 37.077 2.415 37.177 2.515 ;
      RECT 37.077 2.085 37.177 2.185 ;
      RECT 37.077 1.755 37.177 1.855 ;
      RECT 37.077 1.425 37.177 1.525 ;
      RECT 37.077 1.095 37.177 1.195 ;
      RECT 37.077 0.765 37.177 0.865 ;
      RECT 37.223 15.51 37.323 15.61 ;
      RECT 37.223 15.18 37.323 15.28 ;
      RECT 37.223 13.12 37.323 13.22 ;
      RECT 37.223 12.79 37.323 12.89 ;
      RECT 37.302 40.729 37.402 40.829 ;
      RECT 37.302 40.399 37.402 40.499 ;
      RECT 37.302 40.069 37.402 40.169 ;
      RECT 37.302 39.739 37.402 39.839 ;
      RECT 37.302 39.409 37.402 39.509 ;
      RECT 37.302 39.079 37.402 39.179 ;
      RECT 37.302 38.749 37.402 38.849 ;
      RECT 37.302 38.419 37.402 38.519 ;
      RECT 37.302 38.089 37.402 38.189 ;
      RECT 37.302 37.759 37.402 37.859 ;
      RECT 37.302 37.429 37.402 37.529 ;
      RECT 37.302 37.099 37.402 37.199 ;
      RECT 37.302 36.769 37.402 36.869 ;
      RECT 37.302 36.439 37.402 36.539 ;
      RECT 37.407 3.075 37.507 3.175 ;
      RECT 37.407 2.745 37.507 2.845 ;
      RECT 37.407 2.415 37.507 2.515 ;
      RECT 37.407 2.085 37.507 2.185 ;
      RECT 37.407 1.755 37.507 1.855 ;
      RECT 37.407 1.425 37.507 1.525 ;
      RECT 37.407 1.095 37.507 1.195 ;
      RECT 37.407 0.765 37.507 0.865 ;
      RECT 37.553 15.51 37.653 15.61 ;
      RECT 37.553 15.18 37.653 15.28 ;
      RECT 37.553 13.12 37.653 13.22 ;
      RECT 37.553 12.79 37.653 12.89 ;
      RECT 37.632 40.729 37.732 40.829 ;
      RECT 37.632 40.399 37.732 40.499 ;
      RECT 37.632 40.069 37.732 40.169 ;
      RECT 37.632 39.739 37.732 39.839 ;
      RECT 37.632 39.409 37.732 39.509 ;
      RECT 37.632 39.079 37.732 39.179 ;
      RECT 37.632 38.749 37.732 38.849 ;
      RECT 37.632 38.419 37.732 38.519 ;
      RECT 37.632 38.089 37.732 38.189 ;
      RECT 37.632 37.759 37.732 37.859 ;
      RECT 37.632 37.429 37.732 37.529 ;
      RECT 37.632 37.099 37.732 37.199 ;
      RECT 37.632 36.769 37.732 36.869 ;
      RECT 37.632 36.439 37.732 36.539 ;
      RECT 37.737 3.075 37.837 3.175 ;
      RECT 37.737 2.745 37.837 2.845 ;
      RECT 37.737 2.415 37.837 2.515 ;
      RECT 37.737 2.085 37.837 2.185 ;
      RECT 37.737 1.755 37.837 1.855 ;
      RECT 37.737 1.425 37.837 1.525 ;
      RECT 37.737 1.095 37.837 1.195 ;
      RECT 37.737 0.765 37.837 0.865 ;
      RECT 37.883 15.51 37.983 15.61 ;
      RECT 37.883 15.18 37.983 15.28 ;
      RECT 37.883 13.12 37.983 13.22 ;
      RECT 37.883 12.79 37.983 12.89 ;
      RECT 37.962 40.729 38.062 40.829 ;
      RECT 37.962 40.399 38.062 40.499 ;
      RECT 37.962 40.069 38.062 40.169 ;
      RECT 37.962 39.739 38.062 39.839 ;
      RECT 37.962 39.409 38.062 39.509 ;
      RECT 37.962 39.079 38.062 39.179 ;
      RECT 37.962 38.749 38.062 38.849 ;
      RECT 37.962 38.419 38.062 38.519 ;
      RECT 37.962 38.089 38.062 38.189 ;
      RECT 37.962 37.759 38.062 37.859 ;
      RECT 37.962 37.429 38.062 37.529 ;
      RECT 37.962 37.099 38.062 37.199 ;
      RECT 37.962 36.769 38.062 36.869 ;
      RECT 37.962 36.439 38.062 36.539 ;
      RECT 38.067 3.075 38.167 3.175 ;
      RECT 38.067 2.745 38.167 2.845 ;
      RECT 38.067 2.415 38.167 2.515 ;
      RECT 38.067 2.085 38.167 2.185 ;
      RECT 38.067 1.755 38.167 1.855 ;
      RECT 38.067 1.425 38.167 1.525 ;
      RECT 38.067 1.095 38.167 1.195 ;
      RECT 38.067 0.765 38.167 0.865 ;
      RECT 38.213 15.51 38.313 15.61 ;
      RECT 38.213 15.18 38.313 15.28 ;
      RECT 38.213 13.12 38.313 13.22 ;
      RECT 38.213 12.79 38.313 12.89 ;
      RECT 38.292 40.729 38.392 40.829 ;
      RECT 38.292 40.399 38.392 40.499 ;
      RECT 38.292 40.069 38.392 40.169 ;
      RECT 38.292 39.739 38.392 39.839 ;
      RECT 38.292 39.409 38.392 39.509 ;
      RECT 38.292 39.079 38.392 39.179 ;
      RECT 38.292 38.749 38.392 38.849 ;
      RECT 38.292 38.419 38.392 38.519 ;
      RECT 38.292 38.089 38.392 38.189 ;
      RECT 38.292 37.759 38.392 37.859 ;
      RECT 38.292 37.429 38.392 37.529 ;
      RECT 38.292 37.099 38.392 37.199 ;
      RECT 38.292 36.769 38.392 36.869 ;
      RECT 38.292 36.439 38.392 36.539 ;
      RECT 38.397 3.075 38.497 3.175 ;
      RECT 38.397 2.745 38.497 2.845 ;
      RECT 38.397 2.415 38.497 2.515 ;
      RECT 38.397 2.085 38.497 2.185 ;
      RECT 38.397 1.755 38.497 1.855 ;
      RECT 38.397 1.425 38.497 1.525 ;
      RECT 38.397 1.095 38.497 1.195 ;
      RECT 38.397 0.765 38.497 0.865 ;
      RECT 38.543 15.51 38.643 15.61 ;
      RECT 38.543 15.18 38.643 15.28 ;
      RECT 38.543 13.12 38.643 13.22 ;
      RECT 38.543 12.79 38.643 12.89 ;
      RECT 38.622 40.729 38.722 40.829 ;
      RECT 38.622 40.399 38.722 40.499 ;
      RECT 38.622 40.069 38.722 40.169 ;
      RECT 38.622 39.739 38.722 39.839 ;
      RECT 38.622 39.409 38.722 39.509 ;
      RECT 38.622 39.079 38.722 39.179 ;
      RECT 38.622 38.749 38.722 38.849 ;
      RECT 38.622 38.419 38.722 38.519 ;
      RECT 38.622 38.089 38.722 38.189 ;
      RECT 38.622 37.759 38.722 37.859 ;
      RECT 38.622 37.429 38.722 37.529 ;
      RECT 38.622 37.099 38.722 37.199 ;
      RECT 38.622 36.769 38.722 36.869 ;
      RECT 38.622 36.439 38.722 36.539 ;
      RECT 38.727 3.075 38.827 3.175 ;
      RECT 38.727 2.745 38.827 2.845 ;
      RECT 38.727 2.415 38.827 2.515 ;
      RECT 38.727 2.085 38.827 2.185 ;
      RECT 38.727 1.755 38.827 1.855 ;
      RECT 38.727 1.425 38.827 1.525 ;
      RECT 38.727 1.095 38.827 1.195 ;
      RECT 38.727 0.765 38.827 0.865 ;
      RECT 38.873 15.51 38.973 15.61 ;
      RECT 38.873 15.18 38.973 15.28 ;
      RECT 38.873 13.12 38.973 13.22 ;
      RECT 38.873 12.79 38.973 12.89 ;
      RECT 38.952 40.729 39.052 40.829 ;
      RECT 38.952 40.399 39.052 40.499 ;
      RECT 38.952 40.069 39.052 40.169 ;
      RECT 38.952 39.739 39.052 39.839 ;
      RECT 38.952 39.409 39.052 39.509 ;
      RECT 38.952 39.079 39.052 39.179 ;
      RECT 38.952 38.749 39.052 38.849 ;
      RECT 38.952 38.419 39.052 38.519 ;
      RECT 38.952 38.089 39.052 38.189 ;
      RECT 38.952 37.759 39.052 37.859 ;
      RECT 38.952 37.429 39.052 37.529 ;
      RECT 38.952 37.099 39.052 37.199 ;
      RECT 38.952 36.769 39.052 36.869 ;
      RECT 38.952 36.439 39.052 36.539 ;
      RECT 39.203 15.51 39.303 15.61 ;
      RECT 39.203 15.18 39.303 15.28 ;
      RECT 39.203 13.12 39.303 13.22 ;
      RECT 39.203 12.79 39.303 12.89 ;
      RECT 39.282 40.729 39.382 40.829 ;
      RECT 39.282 40.399 39.382 40.499 ;
      RECT 39.282 40.069 39.382 40.169 ;
      RECT 39.282 39.739 39.382 39.839 ;
      RECT 39.282 39.409 39.382 39.509 ;
      RECT 39.282 39.079 39.382 39.179 ;
      RECT 39.282 38.749 39.382 38.849 ;
      RECT 39.282 38.419 39.382 38.519 ;
      RECT 39.282 38.089 39.382 38.189 ;
      RECT 39.282 37.759 39.382 37.859 ;
      RECT 39.282 37.429 39.382 37.529 ;
      RECT 39.282 37.099 39.382 37.199 ;
      RECT 39.282 36.769 39.382 36.869 ;
      RECT 39.282 36.439 39.382 36.539 ;
      RECT 39.533 15.51 39.633 15.61 ;
      RECT 39.533 15.18 39.633 15.28 ;
      RECT 39.533 13.12 39.633 13.22 ;
      RECT 39.533 12.79 39.633 12.89 ;
      RECT 39.612 40.729 39.712 40.829 ;
      RECT 39.612 40.399 39.712 40.499 ;
      RECT 39.612 40.069 39.712 40.169 ;
      RECT 39.612 39.739 39.712 39.839 ;
      RECT 39.612 39.409 39.712 39.509 ;
      RECT 39.612 39.079 39.712 39.179 ;
      RECT 39.612 38.749 39.712 38.849 ;
      RECT 39.612 38.419 39.712 38.519 ;
      RECT 39.612 38.089 39.712 38.189 ;
      RECT 39.612 37.759 39.712 37.859 ;
      RECT 39.612 37.429 39.712 37.529 ;
      RECT 39.612 37.099 39.712 37.199 ;
      RECT 39.612 36.769 39.712 36.869 ;
      RECT 39.612 36.439 39.712 36.539 ;
      RECT 39.863 15.51 39.963 15.61 ;
      RECT 39.863 15.18 39.963 15.28 ;
      RECT 39.863 13.12 39.963 13.22 ;
      RECT 39.863 12.79 39.963 12.89 ;
      RECT 39.942 40.729 40.042 40.829 ;
      RECT 39.942 40.399 40.042 40.499 ;
      RECT 39.942 40.069 40.042 40.169 ;
      RECT 39.942 39.739 40.042 39.839 ;
      RECT 39.942 39.409 40.042 39.509 ;
      RECT 39.942 39.079 40.042 39.179 ;
      RECT 39.942 38.749 40.042 38.849 ;
      RECT 39.942 38.419 40.042 38.519 ;
      RECT 39.942 38.089 40.042 38.189 ;
      RECT 39.942 37.759 40.042 37.859 ;
      RECT 39.942 37.429 40.042 37.529 ;
      RECT 39.942 37.099 40.042 37.199 ;
      RECT 39.942 36.769 40.042 36.869 ;
      RECT 39.942 36.439 40.042 36.539 ;
      RECT 40.193 15.51 40.293 15.61 ;
      RECT 40.193 15.18 40.293 15.28 ;
      RECT 40.193 13.12 40.293 13.22 ;
      RECT 40.193 12.79 40.293 12.89 ;
      RECT 40.272 40.729 40.372 40.829 ;
      RECT 40.272 40.399 40.372 40.499 ;
      RECT 40.272 40.069 40.372 40.169 ;
      RECT 40.272 39.739 40.372 39.839 ;
      RECT 40.272 39.409 40.372 39.509 ;
      RECT 40.272 39.079 40.372 39.179 ;
      RECT 40.272 38.749 40.372 38.849 ;
      RECT 40.272 38.419 40.372 38.519 ;
      RECT 40.272 38.089 40.372 38.189 ;
      RECT 40.272 37.759 40.372 37.859 ;
      RECT 40.272 37.429 40.372 37.529 ;
      RECT 40.272 37.099 40.372 37.199 ;
      RECT 40.272 36.769 40.372 36.869 ;
      RECT 40.272 36.439 40.372 36.539 ;
      RECT 40.523 15.51 40.623 15.61 ;
      RECT 40.523 15.18 40.623 15.28 ;
      RECT 40.523 13.12 40.623 13.22 ;
      RECT 40.523 12.79 40.623 12.89 ;
      RECT 40.602 40.729 40.702 40.829 ;
      RECT 40.602 40.399 40.702 40.499 ;
      RECT 40.602 40.069 40.702 40.169 ;
      RECT 40.602 39.739 40.702 39.839 ;
      RECT 40.602 39.409 40.702 39.509 ;
      RECT 40.602 39.079 40.702 39.179 ;
      RECT 40.602 38.749 40.702 38.849 ;
      RECT 40.602 38.419 40.702 38.519 ;
      RECT 40.602 38.089 40.702 38.189 ;
      RECT 40.602 37.759 40.702 37.859 ;
      RECT 40.602 37.429 40.702 37.529 ;
      RECT 40.602 37.099 40.702 37.199 ;
      RECT 40.602 36.769 40.702 36.869 ;
      RECT 40.602 36.439 40.702 36.539 ;
      RECT 40.853 15.51 40.953 15.61 ;
      RECT 40.853 15.18 40.953 15.28 ;
      RECT 40.853 13.12 40.953 13.22 ;
      RECT 40.853 12.79 40.953 12.89 ;
      RECT 40.932 40.729 41.032 40.829 ;
      RECT 40.932 40.399 41.032 40.499 ;
      RECT 40.932 40.069 41.032 40.169 ;
      RECT 40.932 39.739 41.032 39.839 ;
      RECT 40.932 39.409 41.032 39.509 ;
      RECT 40.932 39.079 41.032 39.179 ;
      RECT 40.932 38.749 41.032 38.849 ;
      RECT 40.932 38.419 41.032 38.519 ;
      RECT 40.932 38.089 41.032 38.189 ;
      RECT 40.932 37.759 41.032 37.859 ;
      RECT 40.932 37.429 41.032 37.529 ;
      RECT 40.932 37.099 41.032 37.199 ;
      RECT 40.932 36.769 41.032 36.869 ;
      RECT 40.932 36.439 41.032 36.539 ;
      RECT 41.183 15.51 41.283 15.61 ;
      RECT 41.183 15.18 41.283 15.28 ;
      RECT 41.183 13.12 41.283 13.22 ;
      RECT 41.183 12.79 41.283 12.89 ;
      RECT 41.262 40.729 41.362 40.829 ;
      RECT 41.262 40.399 41.362 40.499 ;
      RECT 41.262 40.069 41.362 40.169 ;
      RECT 41.262 39.739 41.362 39.839 ;
      RECT 41.262 39.409 41.362 39.509 ;
      RECT 41.262 39.079 41.362 39.179 ;
      RECT 41.262 38.749 41.362 38.849 ;
      RECT 41.262 38.419 41.362 38.519 ;
      RECT 41.262 38.089 41.362 38.189 ;
      RECT 41.262 37.759 41.362 37.859 ;
      RECT 41.262 37.429 41.362 37.529 ;
      RECT 41.262 37.099 41.362 37.199 ;
      RECT 41.262 36.769 41.362 36.869 ;
      RECT 41.262 36.439 41.362 36.539 ;
      RECT 41.513 15.51 41.613 15.61 ;
      RECT 41.513 15.18 41.613 15.28 ;
      RECT 41.513 13.12 41.613 13.22 ;
      RECT 41.513 12.79 41.613 12.89 ;
      RECT 41.592 40.729 41.692 40.829 ;
      RECT 41.592 40.399 41.692 40.499 ;
      RECT 41.592 40.069 41.692 40.169 ;
      RECT 41.592 39.739 41.692 39.839 ;
      RECT 41.592 39.409 41.692 39.509 ;
      RECT 41.592 39.079 41.692 39.179 ;
      RECT 41.592 38.749 41.692 38.849 ;
      RECT 41.592 38.419 41.692 38.519 ;
      RECT 41.592 38.089 41.692 38.189 ;
      RECT 41.592 37.759 41.692 37.859 ;
      RECT 41.592 37.429 41.692 37.529 ;
      RECT 41.592 37.099 41.692 37.199 ;
      RECT 41.592 36.769 41.692 36.869 ;
      RECT 41.592 36.439 41.692 36.539 ;
      RECT 41.843 15.51 41.943 15.61 ;
      RECT 41.843 15.18 41.943 15.28 ;
      RECT 41.843 13.12 41.943 13.22 ;
      RECT 41.843 12.79 41.943 12.89 ;
      RECT 41.922 40.729 42.022 40.829 ;
      RECT 41.922 40.399 42.022 40.499 ;
      RECT 41.922 40.069 42.022 40.169 ;
      RECT 41.922 39.739 42.022 39.839 ;
      RECT 41.922 39.409 42.022 39.509 ;
      RECT 41.922 39.079 42.022 39.179 ;
      RECT 41.922 38.749 42.022 38.849 ;
      RECT 41.922 38.419 42.022 38.519 ;
      RECT 41.922 38.089 42.022 38.189 ;
      RECT 41.922 37.759 42.022 37.859 ;
      RECT 41.922 37.429 42.022 37.529 ;
      RECT 41.922 37.099 42.022 37.199 ;
      RECT 41.922 36.769 42.022 36.869 ;
      RECT 41.922 36.439 42.022 36.539 ;
      RECT 42.173 15.51 42.273 15.61 ;
      RECT 42.173 15.18 42.273 15.28 ;
      RECT 42.173 13.12 42.273 13.22 ;
      RECT 42.173 12.79 42.273 12.89 ;
      RECT 42.252 40.729 42.352 40.829 ;
      RECT 42.252 40.399 42.352 40.499 ;
      RECT 42.252 40.069 42.352 40.169 ;
      RECT 42.252 39.739 42.352 39.839 ;
      RECT 42.252 39.409 42.352 39.509 ;
      RECT 42.252 39.079 42.352 39.179 ;
      RECT 42.252 38.749 42.352 38.849 ;
      RECT 42.252 38.419 42.352 38.519 ;
      RECT 42.252 38.089 42.352 38.189 ;
      RECT 42.252 37.759 42.352 37.859 ;
      RECT 42.252 37.429 42.352 37.529 ;
      RECT 42.252 37.099 42.352 37.199 ;
      RECT 42.252 36.769 42.352 36.869 ;
      RECT 42.252 36.439 42.352 36.539 ;
      RECT 42.503 15.51 42.603 15.61 ;
      RECT 42.503 15.18 42.603 15.28 ;
      RECT 42.503 13.12 42.603 13.22 ;
      RECT 42.503 12.79 42.603 12.89 ;
      RECT 42.582 40.729 42.682 40.829 ;
      RECT 42.582 40.399 42.682 40.499 ;
      RECT 42.582 40.069 42.682 40.169 ;
      RECT 42.582 39.739 42.682 39.839 ;
      RECT 42.582 39.409 42.682 39.509 ;
      RECT 42.582 39.079 42.682 39.179 ;
      RECT 42.582 38.749 42.682 38.849 ;
      RECT 42.582 38.419 42.682 38.519 ;
      RECT 42.582 38.089 42.682 38.189 ;
      RECT 42.582 37.759 42.682 37.859 ;
      RECT 42.582 37.429 42.682 37.529 ;
      RECT 42.582 37.099 42.682 37.199 ;
      RECT 42.582 36.769 42.682 36.869 ;
      RECT 42.582 36.439 42.682 36.539 ;
      RECT 42.912 40.729 43.012 40.829 ;
      RECT 42.912 40.399 43.012 40.499 ;
      RECT 42.912 40.069 43.012 40.169 ;
      RECT 42.912 39.739 43.012 39.839 ;
      RECT 42.912 39.409 43.012 39.509 ;
      RECT 42.912 39.079 43.012 39.179 ;
      RECT 42.912 38.749 43.012 38.849 ;
      RECT 42.912 38.419 43.012 38.519 ;
      RECT 42.912 38.089 43.012 38.189 ;
      RECT 42.912 37.759 43.012 37.859 ;
      RECT 42.912 37.429 43.012 37.529 ;
      RECT 42.912 37.099 43.012 37.199 ;
      RECT 42.912 36.769 43.012 36.869 ;
      RECT 42.912 36.439 43.012 36.539 ;
      RECT 43.242 40.729 43.342 40.829 ;
      RECT 43.242 40.399 43.342 40.499 ;
      RECT 43.242 40.069 43.342 40.169 ;
      RECT 43.242 39.739 43.342 39.839 ;
      RECT 43.242 39.409 43.342 39.509 ;
      RECT 43.242 39.079 43.342 39.179 ;
      RECT 43.242 38.749 43.342 38.849 ;
      RECT 43.242 38.419 43.342 38.519 ;
      RECT 43.242 38.089 43.342 38.189 ;
      RECT 43.242 37.759 43.342 37.859 ;
      RECT 43.242 37.429 43.342 37.529 ;
      RECT 43.242 37.099 43.342 37.199 ;
      RECT 43.242 36.769 43.342 36.869 ;
      RECT 43.242 36.439 43.342 36.539 ;
      RECT 43.572 40.729 43.672 40.829 ;
      RECT 43.572 40.399 43.672 40.499 ;
      RECT 43.572 40.069 43.672 40.169 ;
      RECT 43.572 39.739 43.672 39.839 ;
      RECT 43.572 39.409 43.672 39.509 ;
      RECT 43.572 39.079 43.672 39.179 ;
      RECT 43.572 38.749 43.672 38.849 ;
      RECT 43.572 38.419 43.672 38.519 ;
      RECT 43.572 38.089 43.672 38.189 ;
      RECT 43.572 37.759 43.672 37.859 ;
      RECT 43.572 37.429 43.672 37.529 ;
      RECT 43.572 37.099 43.672 37.199 ;
      RECT 43.572 36.769 43.672 36.869 ;
      RECT 43.572 36.439 43.672 36.539 ;
      RECT 43.902 40.729 44.002 40.829 ;
      RECT 43.902 40.399 44.002 40.499 ;
      RECT 43.902 40.069 44.002 40.169 ;
      RECT 43.902 39.739 44.002 39.839 ;
      RECT 43.902 39.409 44.002 39.509 ;
      RECT 43.902 39.079 44.002 39.179 ;
      RECT 43.902 38.749 44.002 38.849 ;
      RECT 43.902 38.419 44.002 38.519 ;
      RECT 43.902 38.089 44.002 38.189 ;
      RECT 43.902 37.759 44.002 37.859 ;
      RECT 43.902 37.429 44.002 37.529 ;
      RECT 43.902 37.099 44.002 37.199 ;
      RECT 43.902 36.769 44.002 36.869 ;
      RECT 43.902 36.439 44.002 36.539 ;
      RECT 44.232 40.729 44.332 40.829 ;
      RECT 44.232 40.399 44.332 40.499 ;
      RECT 44.232 40.069 44.332 40.169 ;
      RECT 44.232 39.739 44.332 39.839 ;
      RECT 44.232 39.409 44.332 39.509 ;
      RECT 44.232 39.079 44.332 39.179 ;
      RECT 44.232 38.749 44.332 38.849 ;
      RECT 44.232 38.419 44.332 38.519 ;
      RECT 44.232 38.089 44.332 38.189 ;
      RECT 44.232 37.759 44.332 37.859 ;
      RECT 44.232 37.429 44.332 37.529 ;
      RECT 44.232 37.099 44.332 37.199 ;
      RECT 44.232 36.769 44.332 36.869 ;
      RECT 44.232 36.439 44.332 36.539 ;
      RECT 44.383 15.51 44.483 15.61 ;
      RECT 44.383 15.18 44.483 15.28 ;
      RECT 44.383 13.12 44.483 13.22 ;
      RECT 44.383 12.79 44.483 12.89 ;
      RECT 44.562 40.729 44.662 40.829 ;
      RECT 44.562 40.399 44.662 40.499 ;
      RECT 44.562 40.069 44.662 40.169 ;
      RECT 44.562 39.739 44.662 39.839 ;
      RECT 44.562 39.409 44.662 39.509 ;
      RECT 44.562 39.079 44.662 39.179 ;
      RECT 44.562 38.749 44.662 38.849 ;
      RECT 44.562 38.419 44.662 38.519 ;
      RECT 44.562 38.089 44.662 38.189 ;
      RECT 44.562 37.759 44.662 37.859 ;
      RECT 44.562 37.429 44.662 37.529 ;
      RECT 44.562 37.099 44.662 37.199 ;
      RECT 44.562 36.769 44.662 36.869 ;
      RECT 44.562 36.439 44.662 36.539 ;
      RECT 44.713 15.51 44.813 15.61 ;
      RECT 44.713 15.18 44.813 15.28 ;
      RECT 44.713 13.12 44.813 13.22 ;
      RECT 44.713 12.79 44.813 12.89 ;
      RECT 44.892 40.729 44.992 40.829 ;
      RECT 44.892 40.399 44.992 40.499 ;
      RECT 44.892 40.069 44.992 40.169 ;
      RECT 44.892 39.739 44.992 39.839 ;
      RECT 44.892 39.409 44.992 39.509 ;
      RECT 44.892 39.079 44.992 39.179 ;
      RECT 44.892 38.749 44.992 38.849 ;
      RECT 44.892 38.419 44.992 38.519 ;
      RECT 44.892 38.089 44.992 38.189 ;
      RECT 44.892 37.759 44.992 37.859 ;
      RECT 44.892 37.429 44.992 37.529 ;
      RECT 44.892 37.099 44.992 37.199 ;
      RECT 44.892 36.769 44.992 36.869 ;
      RECT 44.892 36.439 44.992 36.539 ;
      RECT 45.043 15.51 45.143 15.61 ;
      RECT 45.043 15.18 45.143 15.28 ;
      RECT 45.043 13.12 45.143 13.22 ;
      RECT 45.043 12.79 45.143 12.89 ;
      RECT 45.222 40.729 45.322 40.829 ;
      RECT 45.222 40.399 45.322 40.499 ;
      RECT 45.222 40.069 45.322 40.169 ;
      RECT 45.222 39.739 45.322 39.839 ;
      RECT 45.222 39.409 45.322 39.509 ;
      RECT 45.222 39.079 45.322 39.179 ;
      RECT 45.222 38.749 45.322 38.849 ;
      RECT 45.222 38.419 45.322 38.519 ;
      RECT 45.222 38.089 45.322 38.189 ;
      RECT 45.222 37.759 45.322 37.859 ;
      RECT 45.222 37.429 45.322 37.529 ;
      RECT 45.222 37.099 45.322 37.199 ;
      RECT 45.222 36.769 45.322 36.869 ;
      RECT 45.222 36.439 45.322 36.539 ;
      RECT 45.373 15.51 45.473 15.61 ;
      RECT 45.373 15.18 45.473 15.28 ;
      RECT 45.373 13.12 45.473 13.22 ;
      RECT 45.373 12.79 45.473 12.89 ;
      RECT 45.552 40.729 45.652 40.829 ;
      RECT 45.552 40.399 45.652 40.499 ;
      RECT 45.552 40.069 45.652 40.169 ;
      RECT 45.552 39.739 45.652 39.839 ;
      RECT 45.552 39.409 45.652 39.509 ;
      RECT 45.552 39.079 45.652 39.179 ;
      RECT 45.552 38.749 45.652 38.849 ;
      RECT 45.552 38.419 45.652 38.519 ;
      RECT 45.552 38.089 45.652 38.189 ;
      RECT 45.552 37.759 45.652 37.859 ;
      RECT 45.552 37.429 45.652 37.529 ;
      RECT 45.552 37.099 45.652 37.199 ;
      RECT 45.552 36.769 45.652 36.869 ;
      RECT 45.552 36.439 45.652 36.539 ;
      RECT 45.703 15.51 45.803 15.61 ;
      RECT 45.703 15.18 45.803 15.28 ;
      RECT 45.703 13.12 45.803 13.22 ;
      RECT 45.703 12.79 45.803 12.89 ;
      RECT 45.882 40.729 45.982 40.829 ;
      RECT 45.882 40.399 45.982 40.499 ;
      RECT 45.882 40.069 45.982 40.169 ;
      RECT 45.882 39.739 45.982 39.839 ;
      RECT 45.882 39.409 45.982 39.509 ;
      RECT 45.882 39.079 45.982 39.179 ;
      RECT 45.882 38.749 45.982 38.849 ;
      RECT 45.882 38.419 45.982 38.519 ;
      RECT 45.882 38.089 45.982 38.189 ;
      RECT 45.882 37.759 45.982 37.859 ;
      RECT 45.882 37.429 45.982 37.529 ;
      RECT 45.882 37.099 45.982 37.199 ;
      RECT 45.882 36.769 45.982 36.869 ;
      RECT 45.882 36.439 45.982 36.539 ;
      RECT 46.033 15.51 46.133 15.61 ;
      RECT 46.033 15.18 46.133 15.28 ;
      RECT 46.033 13.12 46.133 13.22 ;
      RECT 46.033 12.79 46.133 12.89 ;
      RECT 46.212 40.729 46.312 40.829 ;
      RECT 46.212 40.399 46.312 40.499 ;
      RECT 46.212 40.069 46.312 40.169 ;
      RECT 46.212 39.739 46.312 39.839 ;
      RECT 46.212 39.409 46.312 39.509 ;
      RECT 46.212 39.079 46.312 39.179 ;
      RECT 46.212 38.749 46.312 38.849 ;
      RECT 46.212 38.419 46.312 38.519 ;
      RECT 46.212 38.089 46.312 38.189 ;
      RECT 46.212 37.759 46.312 37.859 ;
      RECT 46.212 37.429 46.312 37.529 ;
      RECT 46.212 37.099 46.312 37.199 ;
      RECT 46.212 36.769 46.312 36.869 ;
      RECT 46.212 36.439 46.312 36.539 ;
      RECT 46.363 15.51 46.463 15.61 ;
      RECT 46.363 15.18 46.463 15.28 ;
      RECT 46.363 13.12 46.463 13.22 ;
      RECT 46.363 12.79 46.463 12.89 ;
      RECT 46.542 40.729 46.642 40.829 ;
      RECT 46.542 40.399 46.642 40.499 ;
      RECT 46.542 40.069 46.642 40.169 ;
      RECT 46.542 39.739 46.642 39.839 ;
      RECT 46.542 39.409 46.642 39.509 ;
      RECT 46.542 39.079 46.642 39.179 ;
      RECT 46.542 38.749 46.642 38.849 ;
      RECT 46.542 38.419 46.642 38.519 ;
      RECT 46.542 38.089 46.642 38.189 ;
      RECT 46.542 37.759 46.642 37.859 ;
      RECT 46.542 37.429 46.642 37.529 ;
      RECT 46.542 37.099 46.642 37.199 ;
      RECT 46.542 36.769 46.642 36.869 ;
      RECT 46.542 36.439 46.642 36.539 ;
      RECT 46.693 15.51 46.793 15.61 ;
      RECT 46.693 15.18 46.793 15.28 ;
      RECT 46.693 13.12 46.793 13.22 ;
      RECT 46.693 12.79 46.793 12.89 ;
      RECT 46.872 40.729 46.972 40.829 ;
      RECT 46.872 40.399 46.972 40.499 ;
      RECT 46.872 40.069 46.972 40.169 ;
      RECT 46.872 39.739 46.972 39.839 ;
      RECT 46.872 39.409 46.972 39.509 ;
      RECT 46.872 39.079 46.972 39.179 ;
      RECT 46.872 38.749 46.972 38.849 ;
      RECT 46.872 38.419 46.972 38.519 ;
      RECT 46.872 38.089 46.972 38.189 ;
      RECT 46.872 37.759 46.972 37.859 ;
      RECT 46.872 37.429 46.972 37.529 ;
      RECT 46.872 37.099 46.972 37.199 ;
      RECT 46.872 36.769 46.972 36.869 ;
      RECT 46.872 36.439 46.972 36.539 ;
      RECT 47.023 15.51 47.123 15.61 ;
      RECT 47.023 15.18 47.123 15.28 ;
      RECT 47.023 13.12 47.123 13.22 ;
      RECT 47.023 12.79 47.123 12.89 ;
      RECT 47.202 40.729 47.302 40.829 ;
      RECT 47.202 40.399 47.302 40.499 ;
      RECT 47.202 40.069 47.302 40.169 ;
      RECT 47.202 39.739 47.302 39.839 ;
      RECT 47.202 39.409 47.302 39.509 ;
      RECT 47.202 39.079 47.302 39.179 ;
      RECT 47.202 38.749 47.302 38.849 ;
      RECT 47.202 38.419 47.302 38.519 ;
      RECT 47.202 38.089 47.302 38.189 ;
      RECT 47.202 37.759 47.302 37.859 ;
      RECT 47.202 37.429 47.302 37.529 ;
      RECT 47.202 37.099 47.302 37.199 ;
      RECT 47.202 36.769 47.302 36.869 ;
      RECT 47.202 36.439 47.302 36.539 ;
      RECT 47.353 15.51 47.453 15.61 ;
      RECT 47.353 15.18 47.453 15.28 ;
      RECT 47.353 13.12 47.453 13.22 ;
      RECT 47.353 12.79 47.453 12.89 ;
      RECT 47.532 40.729 47.632 40.829 ;
      RECT 47.532 40.399 47.632 40.499 ;
      RECT 47.532 40.069 47.632 40.169 ;
      RECT 47.532 39.739 47.632 39.839 ;
      RECT 47.532 39.409 47.632 39.509 ;
      RECT 47.532 39.079 47.632 39.179 ;
      RECT 47.532 38.749 47.632 38.849 ;
      RECT 47.532 38.419 47.632 38.519 ;
      RECT 47.532 38.089 47.632 38.189 ;
      RECT 47.532 37.759 47.632 37.859 ;
      RECT 47.532 37.429 47.632 37.529 ;
      RECT 47.532 37.099 47.632 37.199 ;
      RECT 47.532 36.769 47.632 36.869 ;
      RECT 47.532 36.439 47.632 36.539 ;
      RECT 47.683 15.51 47.783 15.61 ;
      RECT 47.683 15.18 47.783 15.28 ;
      RECT 47.683 13.12 47.783 13.22 ;
      RECT 47.683 12.79 47.783 12.89 ;
      RECT 47.862 40.729 47.962 40.829 ;
      RECT 47.862 40.399 47.962 40.499 ;
      RECT 47.862 40.069 47.962 40.169 ;
      RECT 47.862 39.739 47.962 39.839 ;
      RECT 47.862 39.409 47.962 39.509 ;
      RECT 47.862 39.079 47.962 39.179 ;
      RECT 47.862 38.749 47.962 38.849 ;
      RECT 47.862 38.419 47.962 38.519 ;
      RECT 47.862 38.089 47.962 38.189 ;
      RECT 47.862 37.759 47.962 37.859 ;
      RECT 47.862 37.429 47.962 37.529 ;
      RECT 47.862 37.099 47.962 37.199 ;
      RECT 47.862 36.769 47.962 36.869 ;
      RECT 47.862 36.439 47.962 36.539 ;
      RECT 48.013 15.51 48.113 15.61 ;
      RECT 48.013 15.18 48.113 15.28 ;
      RECT 48.013 13.12 48.113 13.22 ;
      RECT 48.013 12.79 48.113 12.89 ;
      RECT 48.192 40.729 48.292 40.829 ;
      RECT 48.192 40.399 48.292 40.499 ;
      RECT 48.192 40.069 48.292 40.169 ;
      RECT 48.192 39.739 48.292 39.839 ;
      RECT 48.192 39.409 48.292 39.509 ;
      RECT 48.192 39.079 48.292 39.179 ;
      RECT 48.192 38.749 48.292 38.849 ;
      RECT 48.192 38.419 48.292 38.519 ;
      RECT 48.192 38.089 48.292 38.189 ;
      RECT 48.192 37.759 48.292 37.859 ;
      RECT 48.192 37.429 48.292 37.529 ;
      RECT 48.192 37.099 48.292 37.199 ;
      RECT 48.192 36.769 48.292 36.869 ;
      RECT 48.192 36.439 48.292 36.539 ;
      RECT 48.343 15.51 48.443 15.61 ;
      RECT 48.343 15.18 48.443 15.28 ;
      RECT 48.343 13.12 48.443 13.22 ;
      RECT 48.343 12.79 48.443 12.89 ;
      RECT 48.522 40.729 48.622 40.829 ;
      RECT 48.522 40.399 48.622 40.499 ;
      RECT 48.522 40.069 48.622 40.169 ;
      RECT 48.522 39.739 48.622 39.839 ;
      RECT 48.522 39.409 48.622 39.509 ;
      RECT 48.522 39.079 48.622 39.179 ;
      RECT 48.522 38.749 48.622 38.849 ;
      RECT 48.522 38.419 48.622 38.519 ;
      RECT 48.522 38.089 48.622 38.189 ;
      RECT 48.522 37.759 48.622 37.859 ;
      RECT 48.522 37.429 48.622 37.529 ;
      RECT 48.522 37.099 48.622 37.199 ;
      RECT 48.522 36.769 48.622 36.869 ;
      RECT 48.522 36.439 48.622 36.539 ;
      RECT 48.673 15.51 48.773 15.61 ;
      RECT 48.673 15.18 48.773 15.28 ;
      RECT 48.673 13.12 48.773 13.22 ;
      RECT 48.673 12.79 48.773 12.89 ;
      RECT 49.003 15.51 49.103 15.61 ;
      RECT 49.003 15.18 49.103 15.28 ;
      RECT 49.003 13.12 49.103 13.22 ;
      RECT 49.003 12.79 49.103 12.89 ;
      RECT 49.333 15.51 49.433 15.61 ;
      RECT 49.333 15.18 49.433 15.28 ;
      RECT 49.333 13.12 49.433 13.22 ;
      RECT 49.333 12.79 49.433 12.89 ;
      RECT 49.663 15.51 49.763 15.61 ;
      RECT 49.663 15.18 49.763 15.28 ;
      RECT 49.663 13.12 49.763 13.22 ;
      RECT 49.663 12.79 49.763 12.89 ;
      RECT 49.993 15.51 50.093 15.61 ;
      RECT 49.993 15.18 50.093 15.28 ;
      RECT 49.993 13.12 50.093 13.22 ;
      RECT 49.993 12.79 50.093 12.89 ;
      RECT 50.323 15.51 50.423 15.61 ;
      RECT 50.323 15.18 50.423 15.28 ;
      RECT 50.323 13.12 50.423 13.22 ;
      RECT 50.323 12.79 50.423 12.89 ;
      RECT 50.653 15.51 50.753 15.61 ;
      RECT 50.653 15.18 50.753 15.28 ;
      RECT 50.653 13.12 50.753 13.22 ;
      RECT 50.653 12.79 50.753 12.89 ;
      RECT 54.26 7.545 54.36 7.645 ;
      RECT 54.26 7.215 54.36 7.315 ;
      RECT 54.26 6.706 54.36 6.806 ;
      RECT 54.26 6.376 54.36 6.476 ;
      RECT 54.59 7.545 54.69 7.645 ;
      RECT 54.59 7.215 54.69 7.315 ;
      RECT 54.59 6.706 54.69 6.806 ;
      RECT 54.59 6.376 54.69 6.476 ;
      RECT 54.92 7.545 55.02 7.645 ;
      RECT 54.92 7.215 55.02 7.315 ;
      RECT 54.92 6.706 55.02 6.806 ;
      RECT 54.92 6.376 55.02 6.476 ;
      RECT 55.25 7.545 55.35 7.645 ;
      RECT 55.25 7.215 55.35 7.315 ;
      RECT 55.25 6.706 55.35 6.806 ;
      RECT 55.25 6.376 55.35 6.476 ;
      RECT 55.58 7.545 55.68 7.645 ;
      RECT 55.58 7.215 55.68 7.315 ;
      RECT 55.58 6.706 55.68 6.806 ;
      RECT 55.58 6.376 55.68 6.476 ;
      RECT 55.91 7.545 56.01 7.645 ;
      RECT 55.91 7.215 56.01 7.315 ;
      RECT 55.91 6.706 56.01 6.806 ;
      RECT 55.91 6.376 56.01 6.476 ;
      RECT 56.829 9.512 56.929 9.612 ;
      RECT 56.829 9.182 56.929 9.282 ;
      RECT 56.829 8.852 56.929 8.952 ;
      RECT 56.829 8.522 56.929 8.622 ;
      RECT 56.829 8.192 56.929 8.292 ;
      RECT 56.829 7.862 56.929 7.962 ;
      RECT 56.829 7.532 56.929 7.632 ;
      RECT 56.829 7.202 56.929 7.302 ;
      RECT 56.829 6.872 56.929 6.972 ;
      RECT 56.829 6.542 56.929 6.642 ;
      RECT 56.829 6.212 56.929 6.312 ;
      RECT 56.829 5.882 56.929 5.982 ;
      RECT 57.159 9.512 57.259 9.612 ;
      RECT 57.159 9.182 57.259 9.282 ;
      RECT 57.159 8.852 57.259 8.952 ;
      RECT 57.159 8.522 57.259 8.622 ;
      RECT 57.159 8.192 57.259 8.292 ;
      RECT 57.159 7.862 57.259 7.962 ;
      RECT 57.159 7.532 57.259 7.632 ;
      RECT 57.159 7.202 57.259 7.302 ;
      RECT 57.159 6.872 57.259 6.972 ;
      RECT 57.159 6.542 57.259 6.642 ;
      RECT 57.159 6.212 57.259 6.312 ;
      RECT 57.159 5.882 57.259 5.982 ;
      RECT 58.139 3.075 58.239 3.175 ;
      RECT 58.139 2.745 58.239 2.845 ;
      RECT 58.139 2.415 58.239 2.515 ;
      RECT 58.139 2.085 58.239 2.185 ;
      RECT 58.139 1.755 58.239 1.855 ;
      RECT 58.139 1.425 58.239 1.525 ;
      RECT 58.139 1.095 58.239 1.195 ;
      RECT 58.139 0.765 58.239 0.865 ;
      RECT 58.469 3.075 58.569 3.175 ;
      RECT 58.469 2.745 58.569 2.845 ;
      RECT 58.469 2.415 58.569 2.515 ;
      RECT 58.469 2.085 58.569 2.185 ;
      RECT 58.469 1.755 58.569 1.855 ;
      RECT 58.469 1.425 58.569 1.525 ;
      RECT 58.469 1.095 58.569 1.195 ;
      RECT 58.469 0.765 58.569 0.865 ;
      RECT 58.799 3.075 58.899 3.175 ;
      RECT 58.799 2.745 58.899 2.845 ;
      RECT 58.799 2.415 58.899 2.515 ;
      RECT 58.799 2.085 58.899 2.185 ;
      RECT 58.799 1.755 58.899 1.855 ;
      RECT 58.799 1.425 58.899 1.525 ;
      RECT 58.799 1.095 58.899 1.195 ;
      RECT 58.799 0.765 58.899 0.865 ;
      RECT 59.129 3.075 59.229 3.175 ;
      RECT 59.129 2.745 59.229 2.845 ;
      RECT 59.129 2.415 59.229 2.515 ;
      RECT 59.129 2.085 59.229 2.185 ;
      RECT 59.129 1.755 59.229 1.855 ;
      RECT 59.129 1.425 59.229 1.525 ;
      RECT 59.129 1.095 59.229 1.195 ;
      RECT 59.129 0.765 59.229 0.865 ;
      RECT 59.459 3.075 59.559 3.175 ;
      RECT 59.459 2.745 59.559 2.845 ;
      RECT 59.459 2.415 59.559 2.515 ;
      RECT 59.459 2.085 59.559 2.185 ;
      RECT 59.459 1.755 59.559 1.855 ;
      RECT 59.459 1.425 59.559 1.525 ;
      RECT 59.459 1.095 59.559 1.195 ;
      RECT 59.459 0.765 59.559 0.865 ;
      RECT 59.789 3.075 59.889 3.175 ;
      RECT 59.789 2.745 59.889 2.845 ;
      RECT 59.789 2.415 59.889 2.515 ;
      RECT 59.789 2.085 59.889 2.185 ;
      RECT 59.789 1.755 59.889 1.855 ;
      RECT 59.789 1.425 59.889 1.525 ;
      RECT 59.789 1.095 59.889 1.195 ;
      RECT 59.789 0.765 59.889 0.865 ;
      RECT 60.119 3.075 60.219 3.175 ;
      RECT 60.119 2.745 60.219 2.845 ;
      RECT 60.119 2.415 60.219 2.515 ;
      RECT 60.119 2.085 60.219 2.185 ;
      RECT 60.119 1.755 60.219 1.855 ;
      RECT 60.119 1.425 60.219 1.525 ;
      RECT 60.119 1.095 60.219 1.195 ;
      RECT 60.119 0.765 60.219 0.865 ;
      RECT 60.449 3.075 60.549 3.175 ;
      RECT 60.449 2.745 60.549 2.845 ;
      RECT 60.449 2.415 60.549 2.515 ;
      RECT 60.449 2.085 60.549 2.185 ;
      RECT 60.449 1.755 60.549 1.855 ;
      RECT 60.449 1.425 60.549 1.525 ;
      RECT 60.449 1.095 60.549 1.195 ;
      RECT 60.449 0.765 60.549 0.865 ;
      RECT 60.779 3.075 60.879 3.175 ;
      RECT 60.779 2.745 60.879 2.845 ;
      RECT 60.779 2.415 60.879 2.515 ;
      RECT 60.779 2.085 60.879 2.185 ;
      RECT 60.779 1.755 60.879 1.855 ;
      RECT 60.779 1.425 60.879 1.525 ;
      RECT 60.779 1.095 60.879 1.195 ;
      RECT 60.779 0.765 60.879 0.865 ;
      RECT 61.109 3.075 61.209 3.175 ;
      RECT 61.109 2.745 61.209 2.845 ;
      RECT 61.109 2.415 61.209 2.515 ;
      RECT 61.109 2.085 61.209 2.185 ;
      RECT 61.109 1.755 61.209 1.855 ;
      RECT 61.109 1.425 61.209 1.525 ;
      RECT 61.109 1.095 61.209 1.195 ;
      RECT 61.109 0.765 61.209 0.865 ;
      RECT 61.439 3.075 61.539 3.175 ;
      RECT 61.439 2.745 61.539 2.845 ;
      RECT 61.439 2.415 61.539 2.515 ;
      RECT 61.439 2.085 61.539 2.185 ;
      RECT 61.439 1.755 61.539 1.855 ;
      RECT 61.439 1.425 61.539 1.525 ;
      RECT 61.439 1.095 61.539 1.195 ;
      RECT 61.439 0.765 61.539 0.865 ;
      RECT 61.769 3.075 61.869 3.175 ;
      RECT 61.769 2.745 61.869 2.845 ;
      RECT 61.769 2.415 61.869 2.515 ;
      RECT 61.769 2.085 61.869 2.185 ;
      RECT 61.769 1.755 61.869 1.855 ;
      RECT 61.769 1.425 61.869 1.525 ;
      RECT 61.769 1.095 61.869 1.195 ;
      RECT 61.769 0.765 61.869 0.865 ;
      RECT 62.099 3.075 62.199 3.175 ;
      RECT 62.099 2.745 62.199 2.845 ;
      RECT 62.099 2.415 62.199 2.515 ;
      RECT 62.099 2.085 62.199 2.185 ;
      RECT 62.099 1.755 62.199 1.855 ;
      RECT 62.099 1.425 62.199 1.525 ;
      RECT 62.099 1.095 62.199 1.195 ;
      RECT 62.099 0.765 62.199 0.865 ;
      RECT 62.429 3.075 62.529 3.175 ;
      RECT 62.429 2.745 62.529 2.845 ;
      RECT 62.429 2.415 62.529 2.515 ;
      RECT 62.429 2.085 62.529 2.185 ;
      RECT 62.429 1.755 62.529 1.855 ;
      RECT 62.429 1.425 62.529 1.525 ;
      RECT 62.429 1.095 62.529 1.195 ;
      RECT 62.429 0.765 62.529 0.865 ;
      RECT 62.759 3.075 62.859 3.175 ;
      RECT 62.759 2.745 62.859 2.845 ;
      RECT 62.759 2.415 62.859 2.515 ;
      RECT 62.759 2.085 62.859 2.185 ;
      RECT 62.759 1.755 62.859 1.855 ;
      RECT 62.759 1.425 62.859 1.525 ;
      RECT 62.759 1.095 62.859 1.195 ;
      RECT 62.759 0.765 62.859 0.865 ;
      RECT 63.089 3.075 63.189 3.175 ;
      RECT 63.089 2.745 63.189 2.845 ;
      RECT 63.089 2.415 63.189 2.515 ;
      RECT 63.089 2.085 63.189 2.185 ;
      RECT 63.089 1.755 63.189 1.855 ;
      RECT 63.089 1.425 63.189 1.525 ;
      RECT 63.089 1.095 63.189 1.195 ;
      RECT 63.089 0.765 63.189 0.865 ;
      RECT 63.419 3.075 63.519 3.175 ;
      RECT 63.419 2.745 63.519 2.845 ;
      RECT 63.419 2.415 63.519 2.515 ;
      RECT 63.419 2.085 63.519 2.185 ;
      RECT 63.419 1.755 63.519 1.855 ;
      RECT 63.419 1.425 63.519 1.525 ;
      RECT 63.419 1.095 63.519 1.195 ;
      RECT 63.419 0.765 63.519 0.865 ;
      RECT 67.475 27.635 67.575 27.735 ;
      RECT 67.475 27.305 67.575 27.405 ;
      RECT 67.475 26.975 67.575 27.075 ;
      RECT 67.475 26.645 67.575 26.745 ;
      RECT 67.475 26.315 67.575 26.415 ;
      RECT 67.475 25.985 67.575 26.085 ;
      RECT 67.475 25.655 67.575 25.755 ;
      RECT 67.475 25.325 67.575 25.425 ;
      RECT 67.475 24.995 67.575 25.095 ;
      RECT 67.475 24.665 67.575 24.765 ;
      RECT 67.475 24.335 67.575 24.435 ;
      RECT 67.475 24.005 67.575 24.105 ;
      RECT 67.475 23.675 67.575 23.775 ;
      RECT 67.475 23.345 67.575 23.445 ;
      RECT 67.805 27.635 67.905 27.735 ;
      RECT 67.805 27.305 67.905 27.405 ;
      RECT 67.805 26.975 67.905 27.075 ;
      RECT 67.805 26.645 67.905 26.745 ;
      RECT 67.805 26.315 67.905 26.415 ;
      RECT 67.805 25.985 67.905 26.085 ;
      RECT 67.805 25.655 67.905 25.755 ;
      RECT 67.805 25.325 67.905 25.425 ;
      RECT 67.805 24.995 67.905 25.095 ;
      RECT 67.805 24.665 67.905 24.765 ;
      RECT 67.805 24.335 67.905 24.435 ;
      RECT 67.805 24.005 67.905 24.105 ;
      RECT 67.805 23.675 67.905 23.775 ;
      RECT 67.805 23.345 67.905 23.445 ;
      RECT 68.135 27.635 68.235 27.735 ;
      RECT 68.135 27.305 68.235 27.405 ;
      RECT 68.135 26.975 68.235 27.075 ;
      RECT 68.135 26.645 68.235 26.745 ;
      RECT 68.135 26.315 68.235 26.415 ;
      RECT 68.135 25.985 68.235 26.085 ;
      RECT 68.135 25.655 68.235 25.755 ;
      RECT 68.135 25.325 68.235 25.425 ;
      RECT 68.135 24.995 68.235 25.095 ;
      RECT 68.135 24.665 68.235 24.765 ;
      RECT 68.135 24.335 68.235 24.435 ;
      RECT 68.135 24.005 68.235 24.105 ;
      RECT 68.135 23.675 68.235 23.775 ;
      RECT 68.135 23.345 68.235 23.445 ;
      RECT 68.465 27.635 68.565 27.735 ;
      RECT 68.465 27.305 68.565 27.405 ;
      RECT 68.465 26.975 68.565 27.075 ;
      RECT 68.465 26.645 68.565 26.745 ;
      RECT 68.465 26.315 68.565 26.415 ;
      RECT 68.465 25.985 68.565 26.085 ;
      RECT 68.465 25.655 68.565 25.755 ;
      RECT 68.465 25.325 68.565 25.425 ;
      RECT 68.465 24.995 68.565 25.095 ;
      RECT 68.465 24.665 68.565 24.765 ;
      RECT 68.465 24.335 68.565 24.435 ;
      RECT 68.465 24.005 68.565 24.105 ;
      RECT 68.465 23.675 68.565 23.775 ;
      RECT 68.465 23.345 68.565 23.445 ;
      RECT 68.795 27.635 68.895 27.735 ;
      RECT 68.795 27.305 68.895 27.405 ;
      RECT 68.795 26.975 68.895 27.075 ;
      RECT 68.795 26.645 68.895 26.745 ;
      RECT 68.795 26.315 68.895 26.415 ;
      RECT 68.795 25.985 68.895 26.085 ;
      RECT 68.795 25.655 68.895 25.755 ;
      RECT 68.795 25.325 68.895 25.425 ;
      RECT 68.795 24.995 68.895 25.095 ;
      RECT 68.795 24.665 68.895 24.765 ;
      RECT 68.795 24.335 68.895 24.435 ;
      RECT 68.795 24.005 68.895 24.105 ;
      RECT 68.795 23.675 68.895 23.775 ;
      RECT 68.795 23.345 68.895 23.445 ;
      RECT 69.125 27.635 69.225 27.735 ;
      RECT 69.125 27.305 69.225 27.405 ;
      RECT 69.125 26.975 69.225 27.075 ;
      RECT 69.125 26.645 69.225 26.745 ;
      RECT 69.125 26.315 69.225 26.415 ;
      RECT 69.125 25.985 69.225 26.085 ;
      RECT 69.125 25.655 69.225 25.755 ;
      RECT 69.125 25.325 69.225 25.425 ;
      RECT 69.125 24.995 69.225 25.095 ;
      RECT 69.125 24.665 69.225 24.765 ;
      RECT 69.125 24.335 69.225 24.435 ;
      RECT 69.125 24.005 69.225 24.105 ;
      RECT 69.125 23.675 69.225 23.775 ;
      RECT 69.125 23.345 69.225 23.445 ;
      RECT 69.455 27.635 69.555 27.735 ;
      RECT 69.455 27.305 69.555 27.405 ;
      RECT 69.455 26.975 69.555 27.075 ;
      RECT 69.455 26.645 69.555 26.745 ;
      RECT 69.455 26.315 69.555 26.415 ;
      RECT 69.455 25.985 69.555 26.085 ;
      RECT 69.455 25.655 69.555 25.755 ;
      RECT 69.455 25.325 69.555 25.425 ;
      RECT 69.455 24.995 69.555 25.095 ;
      RECT 69.455 24.665 69.555 24.765 ;
      RECT 69.455 24.335 69.555 24.435 ;
      RECT 69.455 24.005 69.555 24.105 ;
      RECT 69.455 23.675 69.555 23.775 ;
      RECT 69.455 23.345 69.555 23.445 ;
      RECT 69.785 27.635 69.885 27.735 ;
      RECT 69.785 27.305 69.885 27.405 ;
      RECT 69.785 26.975 69.885 27.075 ;
      RECT 69.785 26.645 69.885 26.745 ;
      RECT 69.785 26.315 69.885 26.415 ;
      RECT 69.785 25.985 69.885 26.085 ;
      RECT 69.785 25.655 69.885 25.755 ;
      RECT 69.785 25.325 69.885 25.425 ;
      RECT 69.785 24.995 69.885 25.095 ;
      RECT 69.785 24.665 69.885 24.765 ;
      RECT 69.785 24.335 69.885 24.435 ;
      RECT 69.785 24.005 69.885 24.105 ;
      RECT 69.785 23.675 69.885 23.775 ;
      RECT 69.785 23.345 69.885 23.445 ;
      RECT 70.115 27.635 70.215 27.735 ;
      RECT 70.115 27.305 70.215 27.405 ;
      RECT 70.115 26.975 70.215 27.075 ;
      RECT 70.115 26.645 70.215 26.745 ;
      RECT 70.115 26.315 70.215 26.415 ;
      RECT 70.115 25.985 70.215 26.085 ;
      RECT 70.115 25.655 70.215 25.755 ;
      RECT 70.115 25.325 70.215 25.425 ;
      RECT 70.115 24.995 70.215 25.095 ;
      RECT 70.115 24.665 70.215 24.765 ;
      RECT 70.115 24.335 70.215 24.435 ;
      RECT 70.115 24.005 70.215 24.105 ;
      RECT 70.115 23.675 70.215 23.775 ;
      RECT 70.115 23.345 70.215 23.445 ;
      RECT 70.445 27.635 70.545 27.735 ;
      RECT 70.445 27.305 70.545 27.405 ;
      RECT 70.445 26.975 70.545 27.075 ;
      RECT 70.445 26.645 70.545 26.745 ;
      RECT 70.445 26.315 70.545 26.415 ;
      RECT 70.445 25.985 70.545 26.085 ;
      RECT 70.445 25.655 70.545 25.755 ;
      RECT 70.445 25.325 70.545 25.425 ;
      RECT 70.445 24.995 70.545 25.095 ;
      RECT 70.445 24.665 70.545 24.765 ;
      RECT 70.445 24.335 70.545 24.435 ;
      RECT 70.445 24.005 70.545 24.105 ;
      RECT 70.445 23.675 70.545 23.775 ;
      RECT 70.445 23.345 70.545 23.445 ;
      RECT 70.775 27.635 70.875 27.735 ;
      RECT 70.775 27.305 70.875 27.405 ;
      RECT 70.775 26.975 70.875 27.075 ;
      RECT 70.775 26.645 70.875 26.745 ;
      RECT 70.775 26.315 70.875 26.415 ;
      RECT 70.775 25.985 70.875 26.085 ;
      RECT 70.775 25.655 70.875 25.755 ;
      RECT 70.775 25.325 70.875 25.425 ;
      RECT 70.775 24.995 70.875 25.095 ;
      RECT 70.775 24.665 70.875 24.765 ;
      RECT 70.775 24.335 70.875 24.435 ;
      RECT 70.775 24.005 70.875 24.105 ;
      RECT 70.775 23.675 70.875 23.775 ;
      RECT 70.775 23.345 70.875 23.445 ;
      RECT 71.105 27.635 71.205 27.735 ;
      RECT 71.105 27.305 71.205 27.405 ;
      RECT 71.105 26.975 71.205 27.075 ;
      RECT 71.105 26.645 71.205 26.745 ;
      RECT 71.105 26.315 71.205 26.415 ;
      RECT 71.105 25.985 71.205 26.085 ;
      RECT 71.105 25.655 71.205 25.755 ;
      RECT 71.105 25.325 71.205 25.425 ;
      RECT 71.105 24.995 71.205 25.095 ;
      RECT 71.105 24.665 71.205 24.765 ;
      RECT 71.105 24.335 71.205 24.435 ;
      RECT 71.105 24.005 71.205 24.105 ;
      RECT 71.105 23.675 71.205 23.775 ;
      RECT 71.105 23.345 71.205 23.445 ;
      RECT 71.435 27.635 71.535 27.735 ;
      RECT 71.435 27.305 71.535 27.405 ;
      RECT 71.435 26.975 71.535 27.075 ;
      RECT 71.435 26.645 71.535 26.745 ;
      RECT 71.435 26.315 71.535 26.415 ;
      RECT 71.435 25.985 71.535 26.085 ;
      RECT 71.435 25.655 71.535 25.755 ;
      RECT 71.435 25.325 71.535 25.425 ;
      RECT 71.435 24.995 71.535 25.095 ;
      RECT 71.435 24.665 71.535 24.765 ;
      RECT 71.435 24.335 71.535 24.435 ;
      RECT 71.435 24.005 71.535 24.105 ;
      RECT 71.435 23.675 71.535 23.775 ;
      RECT 71.435 23.345 71.535 23.445 ;
      RECT 71.765 27.635 71.865 27.735 ;
      RECT 71.765 27.305 71.865 27.405 ;
      RECT 71.765 26.975 71.865 27.075 ;
      RECT 71.765 26.645 71.865 26.745 ;
      RECT 71.765 26.315 71.865 26.415 ;
      RECT 71.765 25.985 71.865 26.085 ;
      RECT 71.765 25.655 71.865 25.755 ;
      RECT 71.765 25.325 71.865 25.425 ;
      RECT 71.765 24.995 71.865 25.095 ;
      RECT 71.765 24.665 71.865 24.765 ;
      RECT 71.765 24.335 71.865 24.435 ;
      RECT 71.765 24.005 71.865 24.105 ;
      RECT 71.765 23.675 71.865 23.775 ;
      RECT 71.765 23.345 71.865 23.445 ;
    LAYER B1 SPACING 0.1 ;
      RECT 41.078 0.72 41.478 3.22 ;
    LAYER B1 ;
      RECT 32.284 13.02 33.124 26.106 ;
      RECT 32.251 13.172 33.158 26.106 ;
      RECT 41.478 0.72 63.655 3.22 ;
  END
  PROPERTY U2DKTabstractName "abstract" ;
END vbbgen_PULPV3_weakdriver

END LIBRARY
