//`define NUM_IF 2 // 4
//`define NUM_OF 2 // 4
`define BANK_SIZE_PARAM 8192
