//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                                      //
// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@8@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@800008@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@88@@@@@@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@@@@@@8CfffffCG8@8CttfC000@@8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@GffttfftffffLLLLC08@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@@@@8Lffff0@@@@@@@@@CftttC800@8@@@@@@@@@@@@@@@@@@@@@@@@@@8LttfftftG@LffG@CfGLLC8@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@@8ffffLCtG@G@8@@@@@@8tf@8t0@08@@@@@@@@@@@@@@@@@@@@@@@@ftttfttfG8LfLCLLffLtC8CfL8@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@GfffffL8@80ftfffC8@@@0GLG@@@@@@@@@@@@@@@@@@@@@@@@@@@@LtttttGtLG0LffGGf0@@8888@@C8@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@8CGLL0@@@@0ttttttttttttttttL@@@8@@@@@@@@@@@@@@@@@@@@@8Lttttt8Ltttt8Lfff0@@@@@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@8C@GG@@@@@@CtttttttttttttttttG@@@@@@@@@@@@@@@@@@@@@@@@8tttL0ftttL@ft@C8@@@@@@@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@0@@@@@8@Ltttttttttttttt1ttf@@@@@@@@@@@@@@@@@@@@@@@@fttfftf8@88@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@@@@@@@@@@@@@@@@8fffttttttt1tttt1ttt10@@@@@@@@@@@@@@@@@@@@@@L11t11ftt8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@@GLC@@@@@@@@@@@0ttC80fttC@@8f1t8LLtttL@@@@@@@@@@@@@@@@@@@@@@8118t0@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@8L8fGGC0@@@@@@@@@CttfftC@8Lft0tt1f0ffC1f@@@@@@@@@@@@@@@@@@@@@@@tt18@@@@@@@@@@@@@@@0CG8@@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@8ffL@@@@@0tf@@@@@Ltttttttttttttt1L111t1f@@@@@@@@@@@@@@@@@@@@@@@@L18@@@@@@@@@@C0@@8@fCGtG@@@@8@@@@@@@@@@@@@ //
// @@@@@@@@@@8000CL@@@088tf@@@GtfC1tttttttt11t101111t@@@@@@@@@@@@@@@@@@@@@@@@@ft@88t8@8@80tttttG8fftfG@@@G@@@@@@@@@@@@@ //
// @@@@@@@@@@@8fG@@@@@@8tft@@@0tf@@@81tt1GG@@@@8t111t@@@@@@@@@@@@@@@@@@@@@@@@@@0fL11f1fGtL80G880ttfffL@fL@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@8G@@@@@@@@@00@@@CL@@@@Gttttttttttt111t@@@@@@@@@@@@@@@@@@@@@@@@@@@@C1tf@8fL@@0@LtL@ffGL88@@@@@@@@@@@@@@@@ //
// @@@@@@@@@@@@CffffC@@@@@@CLG0C08@@@0tfGGf11t1f81t1G@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@1G@t10@@@8LtttLfff@8@@@@@@@@@@@@@@@@ //
// @@@@@@@@LffffftffG0L@@@8fttL@@@@@@801tC@@88@L1f1C@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@0t10@@@@@@@@@Lt8C@@@@@@@@@@@@@@@@@@@ //
// @@@@@@@8fffffffff0080ftL@@@@@@@@@@@@tt1Cf1Ct1ti0@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@0t@@8fC8@Ct@0f@@@@Lf0@@@@@@@@@@@@@@ //
// @@@@@@0ffffL@@@8ffCfLfG@@@@@@@@@@@@@@C1t8L1C1L@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@CG@0ffCttfC@8f8@@@0tL@@@@@@@@@@@@@@ //
// @@@@00CffffffffffC0@@@@@@@@@ttf8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@8@L11fft8@@@@00@@@@8@CtffGf8@@@@@@@@@@@ //
// @@@LffLfCffffffffftf@@@@@@@@tttttf8@@@@@@@08@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ft11t1Ct0f1tttLG08@@0ttffffC@@0tfL8@@@@@@ //
// 8@fG@@@@GffCGGCfffG@@@@@@@@@LtttttttG@@@@GtG@@@@@@@@@@@@@@@@@@@@@@@0GLLCC111tt1t11L010tftttttt@@fffffff0@@@@0fffLfff //
// @L0LLfffLffffffftftL0@@@@@@@@8tttttttt1ttt1@@@@@@@@@@@@@@@@@88i11i111111i1Lt1t@81tt108t0ttttttttfttftfff@@@@@@@CfLff //
// CfffLLfCCC@Cfffftf0tf8@@@@@@@@8ttt1ttt8@811@@@@@@@@@@@@@@@@@i1iC8G11i111GL1t8@@@@0ttttttftttttttf@@Cttff0@@@@@@@@@@@ //
// LLLLLfC8fffLLfffLCL8@@@@@@@@@@@81ttttL@@@Ltf0@@@@@@@@@@@@@@1G@8@80CL1111L8@@tC8tG@@@8CttC@fttLG0@@@CffffC@@@@@@@@@@@ //
// fLLLLf8@ffffffftLff0@@@@@@@@@@@@8tttf0@8fGt11f@@@@@@@@@@@@8tC@@@tL8G1iL8@@@@@t@@88@fttttttttt8@@@@@ffffff@@@@@@@@@@@ //
// 8CffLLGffGGffL08@8@@@@@@Lf@@@@@@@0ttLL@@@ff111@@@@@@@@@@@@@0@Lt8@@t8@8GtfG08G@@@@@G1tttttftttL@@@@@0fffff0@@@@@@@@@@ //
// C@LGL0fLf0@CC@@@8Gff@@@@Lf@@@@@@@@Gttf@@@0111t18@@@@@@@@@@8@f@8@@Gf11ti11111ttttt0Ct080088ftff@@@@@@CffffC@@@@@@@@@@ //
// L@0L00C08@@@0L@@@@@@@@@0f@@@@@@@@@@Ltt@@@81ttttt@@@@@@@@@@@@@@@@@@@@@t1Lt1tttttttttttttttC8@@@@@@@@@LffffL@@@@@@@@@@ //
// @@@@@@@@@@@@@@0C8@@@@8L0@@@@@@@@@@@@ft8@@@8ttCtf@8@@@@@@@@@@@@@@@@@018LtttttttttttttttttttfG@@@@@@@fffffff0@@@@@@@@@ //
// LG@@@@@@@@@@@@@@@@888@@@@@@@@@@@@@@@8t8@@@@LLt0118@@@@@@@@@@@@@@@@@t8CCtttttttttGtLGG0CC008@@@@@@@@CfLffffG@@@@@@@@@ //
// LLC@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@G0@@@@81Gtt0L@@@@@@8@@@@@@@@@@t8@fttLfttttCGtttttffttt8@@@@@@@0ff0fffC@@@@@@@@@ //
// LLG@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@80@@@@@ttfC1L@@@@@@@@@@@@@@@@@t@@tt8@ttttt8GtfG@@000GG@@@@@@@@@ffCfffL@@@@@@@@@ //
// LL8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@C@@@@@L1tt@Gf@@@@@@@@@@@@@@@@8@@tG@@tttCt08ttttttttC@@@@@@@@@@Cffffff8@@@@@@@@ //
// LLLL0@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@L@@@@@8ttt1L@@@@@@@@@@@@@@@@@@@@L8@@8tf@t@@@@8GtLGL0@@@@@@@@@@0ffffff0@@@@@@@@ //
// LLG@@@0G@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@08@@@@@0tttttf@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@LffffLG@@@@@@@@ //
// LLLLG8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@C@@@@@@Lttttt@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@0ffLffL@@@@@@@@ //
// LLC8@@@@@8C@@@@@@@@@@@@@@@@@@@@@@@@@@@@8f8@@@@8ttttt8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@LLLf0f0@@@@@@@ //
// LLLL8@@@0C8@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ff@@@@@8tttC@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@8LL@@CC@@@@@@@ //
//                                                                                                                      //
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Company:        DEI @ UNIBO - University of Bologna                        //
//                                                                            //
// Engineer:       Igor Loi - igor.loi@unibo.it                               //
//                                                                            //
// Additional contributions by:                                               //
//                                                                            //
//                                                                            //
// Create Date:    December 1st 2013                                          //
// Design Name:    Shared instruction cache top module                        //
// Module Name:    icache_top.sv                                              //
// Project Name:   SHARED ICACHE                                              //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    Top module for the Multibank shared instruction cache      //
//                 It supports private configuration, shared with and without //
//                 broadcast capability, and different granularity (1-2-4 WD) //
//                                                                            //
//                                                                            //
// Revision:                                                                  //
// Revision v0.1 - File Created                                               //
// Revision v0.2 - Modified to host the axi based version of the shared $I    //
// Revision v0.3 - Parametric icache                                          //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


`include "ulpsoc_defines.sv"
`include "macro.v"
`timescale 1ns/1ps


module icache_top
#(
    // Parameter for MULTIBANK CACHE
    parameter   NB_CORES                = 4,        // Number of  Processor:     -->  2  |  4  | 8  | 16 | 32
    parameter   NB_REFILL_PORT          = 1,        // DO NOT EDIT --> 1 refill port
    parameter   NB_CACHE_BANKS          = 4,        // Number of  CACHE BANKS:   -->  2  |  4  | 8  | 16 | 32

    parameter   SET_ASSOCIATIVE         = 4,        // 1: DIRECT MAPPED;   2 | 4 | 8    --> Set Associative ICACHE
    parameter   CACHE_LINE              = 1,        // WORDS in each cache line allowed value are 1 - 2 - 4 - 8
    parameter   CACHE_SIZE              = 4096,     // In Byte
    parameter   FIFO_DEPTH              = 2,

    parameter   ICACHE_DATA_WIDTH       = 128,      // 32 | 64 | 128
    parameter   ICACHE_ID_WIDTH         = NB_CORES, // DO NOT EDIT
    parameter   ICACHE_ADDR_WIDTH       = 32,       // DO NOT EDIT

    parameter   L0_BUFFER_FEATURE       = "ENABLED",        // ENABLED | DISABLED
    parameter   L0_SIZE                 = ICACHE_DATA_WIDTH, // DO NOT EDIT

    parameter   INSTR_RDATA_WIDTH       = 32,  // either 32 or ICACHE_DATA_WIDTH

    parameter   SHARED_ICACHE           = "ENABLED",         // ENABLED | DISABLED
    parameter   MULTICAST_FEATURE       = "DISABLED",        // ENABLED | DISABLED
    parameter   MULTICAST_GRANULARITY   = 1,                 // DO NOT EDIT
    parameter   DIRECT_MAPPED_FEATURE   = "DISABLED",         // ENABLED | DISABLED

    parameter   AXI_ID                  = 10,
    parameter   AXI_USER                = 6,
    parameter   AXI_DATA                = 64,
    parameter   AXI_ADDR                = 32
)
(
    // ------------------------------------------------------------------------
    // CORES I$ PLUG ----------------------------------------------------------
    // ------------------------------------------------------------------------
    input logic                                           clk,
    input logic                                           rst_n,
    input logic                                           test_en_i,

    input  logic [NB_CORES-1:0]                           instr_req_i,
    input  logic [NB_CORES-1:0][31:0]                     instr_add_i,
    output logic [NB_CORES-1:0]                           instr_gnt_o,

    output logic [NB_CORES-1:0]                           instr_r_valid_o,
    output logic [NB_CORES-1:0][INSTR_RDATA_WIDTH-1:0]    instr_r_rdata_o,

    // ---------------------------------------------------------------
    // Refill BUS I$ -----------------------------------------
    // ---------------------------------------------------------------
    output logic [AXI_ID-1:0]                             init_awid_o,
    output logic [AXI_ADDR-1:0]                           init_awaddr_o,
    output logic [ 7:0]                                   init_awlen_o,
    output logic [ 2:0]                                   init_awsize_o,
    output logic [ 1:0]                                   init_awburst_o,
    output logic                                          init_awlock_o,
    output logic [ 3:0]                                   init_awcache_o,
    output logic [ 2:0]                                   init_awprot_o,
    output logic [ 3:0]                                   init_awregion_o,
    output logic [ AXI_USER-1:0]                          init_awuser_o,
    output logic [ 3:0]                                   init_awqos_o,
    output logic                                          init_awvalid_o,
    input  logic                                          init_awready_i,

    //AXI write data bus -------------- // // --------------
    output logic  [AXI_DATA-1:0]                          init_wdata_o,
    output logic  [AXI_DATA/8-1:0]                        init_wstrb_o,
    output logic                                          init_wlast_o,
    output logic  [ AXI_USER-1:0]                         init_wuser_o,
    output logic                                          init_wvalid_o,
    input  logic                                          init_wready_i,
    // ---------------------------------------------------------------

    //AXI BACKWARD write response bus -------------- // // --------------
    input  logic  [AXI_ID-1:0]                            init_bid_i,
    input  logic  [ 1:0]                                  init_bresp_i,
    input  logic  [ AXI_USER-1:0]                         init_buser_i,
    input  logic                                          init_bvalid_i,
    output logic                                          init_bready_o,
    // ---------------------------------------------------------------

    //AXI read address bus -------------------------------------------
    output  logic [AXI_ID-1:0]                            init_arid_o,       //
    output  logic [AXI_ADDR-1:0]                          init_araddr_o,     //
    output  logic [ 7:0]                                  init_arlen_o,      // burst length - 1 to 256
    output  logic [ 2:0]                                  init_arsize_o,     // size of each transfer in burst
    output  logic [ 1:0]                                  init_arburst_o,    // for bursts>1, accept only incr burst=01
    output  logic                                         init_arlock_o,     // only normal access supported axs_awlock=00
    output  logic [ 3:0]                                  init_arcache_o,    //
    output  logic [ 2:0]                                  init_arprot_o,     //
    output  logic [ 3:0]                                  init_arregion_o,   //
    output  logic [ AXI_USER-1:0]                         init_aruser_o,     //
    output  logic [ 3:0]                                  init_arqos_o,      //
    output  logic                                         init_arvalid_o,    // master addr valid
    input logic                                           init_arready_i,    // slave ready to accept
    // --------------------------------------------------------------------------------

    //AXI BACKWARD read data bus ----------------------------------------------
    input  logic [AXI_ID-1:0]                             init_rid_i,        //
    input  logic [AXI_DATA-1:0]                           init_rdata_i,      //
    input  logic [ 1:0]                                   init_rresp_i,      //
    input  logic                                          init_rlast_i,      // last transfer in burst
    input  logic [ AXI_USER-1:0]                          init_ruser_i,      //
    input  logic                                          init_rvalid_i,     // slave data valid
    output logic                                          init_rready_o,     // master ready to accept
    // Control ports
    ICACHE_CTRL_UNIT_BUS.Slave                            IC_ctrl_unit_slave_if[NB_CACHE_BANKS],
    L0_CTRL_UNIT_BUS.Slave                                L0_ctrl_unit_slave_if[NB_CORES]
);


   localparam  OFFSET_BIT  =  2;
   localparam  BLI_LSB     =  OFFSET_BIT  + `log2(CACHE_LINE-1);
   localparam  BLI_MSB     =  OFFSET_BIT  + `log2(CACHE_LINE-1)+`log2(NB_CACHE_BANKS-1)-1;
   localparam  AXI_ID_INT  =  1;
   localparam  AXI_ID_OUT  =  `log2(NB_CACHE_BANKS-1) + 1;
   genvar      i,k,j,w,z;


   logic icache_is_private;

   assign icache_is_private = IC_ctrl_unit_slave_if[0].icache_is_private;



  // AXI BUSSES BETWEEN CACHE BANKS and AXI NODE
  //AXI write address bus -------------- // // --------------
  logic [NB_CACHE_BANKS-1:0][AXI_ID_INT-1:0]                 init_awid_internal;       //
  logic [NB_CACHE_BANKS-1:0][AXI_ADDR-1:0]                   init_awaddr_internal;     //
  logic [NB_CACHE_BANKS-1:0][ 7:0]                           init_awlen_internal;      // burst length 0-255 beat
  logic [NB_CACHE_BANKS-1:0][ 2:0]                           init_awsize_internal;     // size of each transfer in burst
  logic [NB_CACHE_BANKS-1:0][ 1:0]                           init_awburst_internal;    // for bursts>1; accept only incr burst=01
  logic [NB_CACHE_BANKS-1:0]                                 init_awlock_internal;     // only normal access supported axs_awlock=00
  logic [NB_CACHE_BANKS-1:0][ 3:0]                           init_awcache_internal;    //
  logic [NB_CACHE_BANKS-1:0][ 2:0]                           init_awprot_internal;     //
  logic [NB_CACHE_BANKS-1:0][ 3:0]                           init_awregion_internal;   //
  logic [NB_CACHE_BANKS-1:0][ AXI_USER-1:0]                  init_awuser_internal;     //
  logic [NB_CACHE_BANKS-1:0][ 3:0]                           init_awqos_internal;      //
  logic [NB_CACHE_BANKS-1:0]                                 init_awvalid_internal;    // master addr valid
  logic [NB_CACHE_BANKS-1:0]                                 init_awready_internal;    // slave ready to accept
  // ---------------------------------------------------------------

  //AXI write data bus -------------- // // --------------
  logic [NB_CACHE_BANKS-1:0] [AXI_DATA-1:0]                  init_wdata_internal;
  logic [NB_CACHE_BANKS-1:0] [AXI_DATA/8-1:0]                init_wstrb_internal;      // 1 strobe per byte
  logic [NB_CACHE_BANKS-1:0]                                 init_wlast_internal;      // last transfer in burst
  logic [NB_CACHE_BANKS-1:0] [ AXI_USER-1:0]                 init_wuser_internal;      // user sideband signals
  logic [NB_CACHE_BANKS-1:0]                                 init_wvalid_internal;     // master data valid
  logic [NB_CACHE_BANKS-1:0]                                 init_wready_internal;     // slave ready to accept
  // ---------------------------------------------------------------

  //AXI BACKWARD write response bus -------------- // // --------------
  logic [NB_CACHE_BANKS-1:0] [AXI_ID_INT-1:0]                init_bid_internal;
  logic [NB_CACHE_BANKS-1:0] [ 1:0]                          init_bresp_internal;
  logic [NB_CACHE_BANKS-1:0] [ AXI_USER-1:0]                 init_buser_internal;
  logic [NB_CACHE_BANKS-1:0]                                 init_bvalid_internal;
  logic [NB_CACHE_BANKS-1:0]                                 init_bready_internal;
  // ---------------------------------------------------------------

  //AXI read address bus -------------------------------------------
  logic [NB_CACHE_BANKS-1:0][AXI_ID_INT-1:0]                 init_arid_internal;
  logic [NB_CACHE_BANKS-1:0][AXI_ADDR-1:0]                   init_araddr_internal;
  logic [NB_CACHE_BANKS-1:0][ 7:0]                           init_arlen_internal;      // burst length - 1 to 16
  logic [NB_CACHE_BANKS-1:0][ 2:0]                           init_arsize_internal;     // size of each transfer in burst
  logic [NB_CACHE_BANKS-1:0][ 1:0]                           init_arburst_internal;    // for bursts>1; accept only incr burst=01
  logic [NB_CACHE_BANKS-1:0]                                 init_arlock_internal;     // only normal access supported axs_awlock=00
  logic [NB_CACHE_BANKS-1:0][ 3:0]                           init_arcache_internal;    //
  logic [NB_CACHE_BANKS-1:0][ 2:0]                           init_arprot_internal;     //
  logic [NB_CACHE_BANKS-1:0][ 3:0]                           init_arregion_internal;   //
  logic [NB_CACHE_BANKS-1:0][ AXI_USER-1:0]                  init_aruser_internal;     //
  logic [NB_CACHE_BANKS-1:0][ 3:0]                           init_arqos_internal;      //
  logic [NB_CACHE_BANKS-1:0]                                 init_arvalid_internal;    // master addr valid
  logic [NB_CACHE_BANKS-1:0]                                 init_arready_internal;    // slave ready to accept
  // ---------------------------------------------------------------

  //AXI BACKWARD read data bus ----------------------------------------------
  logic [NB_CACHE_BANKS-1:0][AXI_ID_INT-1:0]                 init_rid_internal;     //
  logic [NB_CACHE_BANKS-1:0][AXI_DATA-1:0]                   init_rdata_internal;   //
  logic [NB_CACHE_BANKS-1:0][ 1:0]                           init_rresp_internal;   //
  logic [NB_CACHE_BANKS-1:0]                                 init_rlast_internal;   // last transfer in burst
  logic [NB_CACHE_BANKS-1:0][AXI_USER-1:0]                   init_ruser_internal;   //
  logic [NB_CACHE_BANKS-1:0]                                 init_rvalid_internal;  // slave data valid
  logic [NB_CACHE_BANKS-1:0]                                 init_rready_internal;  // master ready to accept



  // Signal From Fetch Buffer to Shared icache Interconnect
  logic [NB_CORES-1:0]                                       instr_req_FB_to_IC;
  logic [NB_CORES-1:0][ICACHE_ADDR_WIDTH-1:0]                instr_add_FB_to_IC;
  logic [NB_CORES-1:0]                                       instr_gnt_FB_to_IC;
  logic [NB_CORES-1:0]                                       instr_r_valid_FB_to_IC;
  logic [NB_CORES-1:0][ICACHE_DATA_WIDTH-1:0]                instr_r_rdata_FB_to_IC;


////////////////////////////////////////////////////////////
// ██╗      ██████╗     ██████╗ ██╗   ██╗███████╗███████╗ //
// ██║     ██╔═████╗    ██╔══██╗██║   ██║██╔════╝██╔════╝ //
// ██║     ██║██╔██║    ██████╔╝██║   ██║█████╗  █████╗   //
// ██║     ████╔╝██║    ██╔══██╗██║   ██║██╔══╝  ██╔══╝   //
// ███████╗╚██████╔╝    ██████╔╝╚██████╔╝██║     ██║      //
// ╚══════╝ ╚═════╝     ╚═════╝  ╚═════╝ ╚═╝     ╚═╝      //
////////////////////////////////////////////////////////////
generate

for (k=0;k<NB_CORES;k++)
begin : FETCH_BUFFER
    if(L0_BUFFER_FEATURE == "ENABLED")
    begin : _L0_ENABLED_

          case(L0_SIZE)
          32:
          begin : _32_BIT_
                fetch_buffer_32 fetch_buffer_i
                (
                    .clk              (  clk                       ),
                    .rst_n            (  rst_n                     ),

                    .instr_req_i      (  instr_req_i[k]            ),
                    .instr_add_i      (  instr_add_i[k]            ),
                    .instr_gnt_o      (  instr_gnt_o[k]            ),

                    .instr_r_valid_o  (  instr_r_valid_o[k]        ),
                    .instr_r_rdata_o  (  instr_r_rdata_o[k]        ),

                    .instr_req_o      (  instr_req_FB_to_IC[k]     ),
                    .instr_add_o      (  instr_add_FB_to_IC[k]     ),
                    .instr_gnt_i      (  instr_gnt_FB_to_IC[k]     ),

                    .instr_r_valid_i  (  instr_r_valid_FB_to_IC[k] ),
                    .instr_r_rdata_i  (  instr_r_rdata_FB_to_IC[k] )
                );
          end

          64:
          begin : _64_BIT_
                fetch_buffer_64 fetch_buffer_i
                (
                    .clk              (  clk                       ),
                    .rst_n            (  rst_n                     ),

                    .instr_req_i      (  instr_req_i[k]            ),
                    .instr_add_i      (  instr_add_i[k]            ),
                    .instr_gnt_o      (  instr_gnt_o[k]            ),

                    .instr_r_valid_o  (  instr_r_valid_o[k]        ),
                    .instr_r_rdata_o  (  instr_r_rdata_o[k]        ),

                    .instr_req_o      (  instr_req_FB_to_IC[k]     ),
                    .instr_add_o      (  instr_add_FB_to_IC[k]     ),
                    .instr_gnt_i      (  instr_gnt_FB_to_IC[k]     ),

                    .instr_r_valid_i  (  instr_r_valid_FB_to_IC[k] ),
                    .instr_r_rdata_i  (  instr_r_rdata_FB_to_IC[k] )
                );
          end

          128:
          begin : _128_BIT_
                fetch_buffer_128 fetch_buffer_i
                (
                    .flush_i          (  L0_ctrl_unit_slave_if[k].flush_FetchBuffer    ),
                    .ack_flush_o      (  L0_ctrl_unit_slave_if[k].flush_ack            ),
                    .clk              (  clk                       ),
                    .rst_n            (  rst_n                     ),

                    .instr_req_i      (  instr_req_i[k]            ),
                    .instr_add_i      (  instr_add_i[k]            ),
                    .instr_gnt_o      (  instr_gnt_o[k]            ),

                    .instr_r_valid_o  (  instr_r_valid_o[k]        ),
                    .instr_r_rdata_o  (  instr_r_rdata_o[k]        ),


                    .instr_req_o      (  instr_req_FB_to_IC[k]     ),
                    .instr_add_o      (  instr_add_FB_to_IC[k]     ),
                    .instr_gnt_i      (  instr_gnt_FB_to_IC[k]     ),

                    .instr_r_valid_i  (  instr_r_valid_FB_to_IC[k] ),
                    .instr_r_rdata_i  (  instr_r_rdata_FB_to_IC[k] )
                );
          end


          // REMOVE THE FETCH BUFFER
          default :
          begin : _OUT_OF_RANGE_
                assign instr_r_valid_o[k]     = instr_r_valid_FB_to_IC[k];
                assign instr_r_rdata_o[k]     = instr_r_rdata_FB_to_IC[k];
                assign instr_gnt_o[k]         = instr_gnt_FB_to_IC[k];
                assign instr_req_FB_to_IC[k]  = instr_req_i[k];
                assign instr_add_FB_to_IC[k]  = instr_add_i[k];
          end

          endcase

  end
  else //else (L0_BUFFER_FEATURE == "ENABLED")
  begin : _NO_L0_BUFFER_
          assign instr_r_valid_o[k]                = instr_r_valid_FB_to_IC[k];
          assign instr_r_rdata_o[k]                = instr_r_rdata_FB_to_IC[k];
          assign instr_gnt_o[k]                    = instr_gnt_FB_to_IC[k];
          assign instr_req_FB_to_IC[k]             = instr_req_i[k];
          assign instr_add_FB_to_IC[k]             = instr_add_i[k];
  end
end
endgenerate



///////////////////////////////////////////////////////////////////////////////////////////
// ██╗ ██████╗ █████╗  ██████╗██╗  ██╗███████╗        ██████╗  █████╗ ███╗   ██╗██╗  ██╗ //
// ██║██╔════╝██╔══██╗██╔════╝██║  ██║██╔════╝        ██╔══██╗██╔══██╗████╗  ██║██║ ██╔╝ //
// ██║██║     ███████║██║     ███████║█████╗          ██████╔╝███████║██╔██╗ ██║█████╔╝  //
// ██║██║     ██╔══██║██║     ██╔══██║██╔══╝          ██╔══██╗██╔══██║██║╚██╗██║██╔═██╗  //
// ██║╚██████╗██║  ██║╚██████╗██║  ██║███████╗███████╗██████╔╝██║  ██║██║ ╚████║██║  ██╗ //
// ╚═╝ ╚═════╝╚═╝  ╚═╝ ╚═════╝╚═╝  ╚═╝╚══════╝╚══════╝╚═════╝ ╚═╝  ╚═╝╚═╝  ╚═══╝╚═╝  ╚═╝ //
///////////////////////////////////////////////////////////////////////////////////////////
generate

if(SHARED_ICACHE == "ENABLED")
begin : _SHARED_ENABLED_
   // -------------------------------------------------------------------------
   // SHARED_ICACHE_INTERCONNECT (intc) to ICACHE BANKS  (cb) signals ---------
   // -------------------------------------------------------------------------
   logic [NB_CACHE_BANKS-1:0]                                  fetch_req_intc_to_cb;
   logic [NB_CACHE_BANKS-1:0]                                  fetch_grant_cb_to_intc;
   logic [NB_CACHE_BANKS-1:0][ICACHE_ADDR_WIDTH-1:0]           fetch_addr_intc_to_cb;
   logic [NB_CACHE_BANKS-1:0][ICACHE_ID_WIDTH-1:0]             fetch_ID_intc_to_cb;

   logic [NB_CACHE_BANKS-1:0][ICACHE_DATA_WIDTH-1:0]           fetch_r_rdata_cb_to_intc;
   logic [NB_CACHE_BANKS-1:0]                                  fetch_r_valid_cb_to_intc;
   logic [NB_CACHE_BANKS-1:0][ICACHE_ID_WIDTH-1:0]             fetch_r_ID_cb_to_intc;

   // -------------------------------------------------------------------------
   // SHARED_ICACHE_INTERCONNECT                                      ---------
   // -------------------------------------------------------------------------
   XBAR_ICACHE
   #(
       .N_CH0                 ( NB_CORES                                                                             ),  //--> CH0
       .N_CH1                 ( 0                                                                                    ),  //--> CH1 , not used
       .N_SLAVE               ( NB_CACHE_BANKS                                                                       ),
       .BLI_LSB               ( OFFSET_BIT + `log2((ICACHE_DATA_WIDTH/32)*CACHE_LINE-1)                              ),
       .BLI_MSB               ( OFFSET_BIT + `log2((ICACHE_DATA_WIDTH/32)*CACHE_LINE-1) + `log2(NB_CACHE_BANKS-1) -1 ),
       .MULTICAST_FEATURE     ( MULTICAST_FEATURE                                                                    ),
       .MULTICAST_GRANULARITY ( MULTICAST_GRANULARITY                                                                ),
       .ADDR_WIDTH            ( ICACHE_ADDR_WIDTH                                                                    ),
       .DATA_WIDTH            ( ICACHE_DATA_WIDTH                                                                    )
   )
   ICACHE_INTERCONNECT
   (
      // ---------------- Cores Side   -----------------------------------------------------------
      .data_req_i          (   instr_req_FB_to_IC       ),            // Data request
      .data_add_i          (   instr_add_FB_to_IC       ),            // Data request Address
      .data_gnt_o          (   instr_gnt_FB_to_IC       ),        // Grant Incoming Request

      .data_r_valid_o      (   instr_r_valid_FB_to_IC   ),            // Data Response Valid (For LOAD/STORE commands)
      .data_r_rdata_o      (   instr_r_rdata_FB_to_IC   ),             // Data Response DATA (For LOAD commands)

      // ---------------- ICACHE BANKS SIDE (Interleaving--> Cache Line) --------------------------
      .data_req_o          (   fetch_req_intc_to_cb     ),         // Data request
      .data_add_o          (   fetch_addr_intc_to_cb    ),         // Data request Address
      .data_ID_o           (   fetch_ID_intc_to_cb      ),         // Data request Address
      .data_gnt_i          (   fetch_grant_cb_to_intc   ),             // Data Grant

      .data_r_valid_i      (   fetch_r_valid_cb_to_intc ),            // valid REspone (must be accepted always)
      .data_r_ID_i         (   fetch_r_ID_cb_to_intc    ),             // Data Response ID (For LOAD commands)
      .data_r_rdata_i      (   fetch_r_rdata_cb_to_intc ),             // Data Response DATA (For LOAD and STORE)

      .clk                 (   clk                      ),
      .rst_n               (   rst_n                    ),
      .icache_is_private_i (   icache_is_private        )
   );




   // -------------------------------------------------------------------------
   // SHARED_ICACHE BANKS                                             ---------
   // -------------------------------------------------------------------------
   for(i=0; i<NB_CACHE_BANKS; i++)
   begin : SHARED_ICACHE_BANKS
         icache
         #(
            .N_BANKS                ( NB_CACHE_BANKS                 ),
            .SET_ASSOCIATIVE        ( SET_ASSOCIATIVE                ),
            .CACHE_LINE             ( CACHE_LINE                     ),
            .CACHE_SIZE             ( CACHE_SIZE/NB_CACHE_BANKS      ),  //In Byte
            .CACHE_ID               ( i                              ),
            .FIFO_DEPTH             ( FIFO_DEPTH                     ),

            .ICACHE_DATA_WIDTH      ( ICACHE_DATA_WIDTH              ),
            .ICACHE_ID_WIDTH        ( ICACHE_ID_WIDTH                ),
            .ICACHE_ADDR_WIDTH      ( ICACHE_ADDR_WIDTH              ),

            .DIRECT_MAPPED_FEATURE  ( DIRECT_MAPPED_FEATURE          ),

            .AXI_ID                 ( AXI_ID_INT                     ),
            .AXI_ADDR               ( AXI_ADDR                       ),
            .AXI_DATA               ( AXI_DATA                       ),
            .AXI_USER               ( AXI_USER                       )
         )
         u_icache_bank
         (
            // ---------------------------------------------------------------
            // I/O Port Declarations -----------------------------------------
            // ---------------------------------------------------------------
            .clk             ( clk                            ),
            .rst_n           ( rst_n                          ),
            .test_en_i       ( test_en_i                      ),
            .icache_is_private_i ( icache_is_private          ),

            // ---------------------------------------------------------------
            // SHARED_ICACHE_INTERCONNECT Port Declarations -----------------------------------------
            // ---------------------------------------------------------------
            .fetch_req_i     (  fetch_req_intc_to_cb[i]      ),
            .fetch_grant_o   (  fetch_grant_cb_to_intc[i]    ),
            .fetch_addr_i    (  fetch_addr_intc_to_cb[i]     ),
            .fetch_ID_i      (  fetch_ID_intc_to_cb[i]       ),
            .fetch_r_rdata_o (  fetch_r_rdata_cb_to_intc[i]  ),
            .fetch_r_valid_o (  fetch_r_valid_cb_to_intc[i]  ),
            .fetch_r_ID_o    (  fetch_r_ID_cb_to_intc[i]     ),

            // §§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§ //
            // §§§§§§§§§§§§§§§§§§§    REFILL Request side  §§§§§§§§§§§§§§§§§§§§§§§ //
            // §§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§ //
            .init_awid_o     (  init_awid_internal[i]     ),
            .init_awaddr_o   (  init_awaddr_internal[i]   ),
            .init_awlen_o    (  init_awlen_internal[i]    ),
            .init_awsize_o   (  init_awsize_internal[i]   ),
            .init_awburst_o  (  init_awburst_internal[i]  ),
            .init_awlock_o   (  init_awlock_internal[i]   ),
            .init_awcache_o  (  init_awcache_internal[i]  ),
            .init_awprot_o   (  init_awprot_internal[i]   ),
            .init_awregion_o (  init_awregion_internal[i] ),
            .init_awuser_o   (  init_awuser_internal[i]   ),
            .init_awqos_o    (  init_awqos_internal[i]    ),
            .init_awvalid_o  (  init_awvalid_internal[i]  ),
            .init_awready_i  (  init_awready_internal[i]  ),

            .init_wdata_o    (  init_wdata_internal[i]    ),
            .init_wstrb_o    (  init_wstrb_internal[i]    ),
            .init_wlast_o    (  init_wlast_internal[i]    ),
            .init_wuser_o    (  init_wuser_internal[i]    ),
            .init_wvalid_o   (  init_wvalid_internal[i]   ),
            .init_wready_i   (  init_wready_internal[i]   ),

            .init_bid_i      (  init_bid_internal[i]      ),
            .init_bresp_i    (  init_bresp_internal[i]    ),
            .init_buser_i    (  init_buser_internal[i]    ),
            .init_bvalid_i   (  init_bvalid_internal[i]   ),
            .init_bready_o   (  init_bready_internal[i]   ),

            .init_arid_o     (  init_arid_internal[i]     ),
            .init_araddr_o   (  init_araddr_internal[i]   ),
            .init_arlen_o    (  init_arlen_internal[i]    ),
            .init_arsize_o   (  init_arsize_internal[i]   ),
            .init_arburst_o  (  init_arburst_internal[i]  ),
            .init_arlock_o   (  init_arlock_internal[i]   ),
            .init_arcache_o  (  init_arcache_internal[i]  ),
            .init_arprot_o   (  init_arprot_internal[i]   ),
            .init_arregion_o (  init_arregion_internal[i] ),
            .init_aruser_o   (  init_aruser_internal[i]   ),
            .init_arqos_o    (  init_arqos_internal[i]    ),
            .init_arvalid_o  (  init_arvalid_internal[i]  ),
            .init_arready_i  (  init_arready_internal[i]  ),

            .init_rid_i     (  init_rid_internal[i]       ),
            .init_rdata_i   (  init_rdata_internal[i]     ),
            .init_rresp_i   (  init_rresp_internal[i]     ),
            .init_rlast_i   (  init_rlast_internal[i]     ),
            .init_ruser_i   (  init_ruser_internal[i]     ),
            .init_rvalid_i  (  init_rvalid_internal[i]    ),
            .init_rready_o  (  init_rready_internal[i]    ),

            // Control ports
            .ctrl_req_enable_icache_i      ( IC_ctrl_unit_slave_if[i].ctrl_req_enable    ),
            .ctrl_ack_enable_icache_o      ( IC_ctrl_unit_slave_if[i].ctrl_ack_enable    ),
            .ctrl_req_disable_icache_i     ( IC_ctrl_unit_slave_if[i].ctrl_req_disable   ),
            .ctrl_ack_disable_icache_o     ( IC_ctrl_unit_slave_if[i].ctrl_ack_disable   ),
            .ctrl_pending_trans_icache_o   ( IC_ctrl_unit_slave_if[i].ctrl_pending_trans )
`ifdef FEATURE_ICACHE_STAT
            ,
            .ctrl_hit_count_icache_o       ( IC_ctrl_unit_slave_if[i].ctrl_hit_count     ),
            .ctrl_trans_count_icache_o     ( IC_ctrl_unit_slave_if[i].ctrl_trans_count   ),
            .ctrl_clear_regs_icache_i      ( IC_ctrl_unit_slave_if[i].ctrl_clear_regs    ),
            .ctrl_enable_regs_icache_i     ( IC_ctrl_unit_slave_if[i].ctrl_enable_regs   )
`endif
         );
   end // ~for(i=0; i<NB_CACHE_BANKS; i++) --> inst icache_bank
end // ~if(SHARED_ICACHE == "ENABLED")
else //  PRIVATE ICACHE BANKS
begin : GEN_PRI
            for(i=0; i<NB_CORES; i++)
            begin : PRIVATE_ICACHE_BANKS
              icache
              #(
                  .N_BANKS                 ( 1                      ),
                  .SET_ASSOCIATIVE         ( SET_ASSOCIATIVE        ),
                  .CACHE_LINE              ( CACHE_LINE             ),
                  .CACHE_SIZE              ( CACHE_SIZE             ),  //In Byte
                  .CACHE_ID                ( i                      ),
                  .FIFO_DEPTH              ( FIFO_DEPTH             ),

                  .ICACHE_DATA_WIDTH       ( ICACHE_DATA_WIDTH      ),
                  .ICACHE_ID_WIDTH         ( ICACHE_ID_WIDTH        ),
                  .ICACHE_ADDR_WIDTH       ( ICACHE_ADDR_WIDTH      ),

                  .DIRECT_MAPPED_FEATURE   ( DIRECT_MAPPED_FEATURE  ),

                  .AXI_ID                  ( AXI_ID_INT             ),
                  .AXI_ADDR                ( AXI_ADDR               ),
                  .AXI_DATA                ( AXI_DATA               ),
                  .AXI_USER                ( AXI_USER               )
              )
              u_icache_bank
              (
                  // ---------------------------------------------------------------
                  // I/O Port Declarations -----------------------------------------
                  // ---------------------------------------------------------------
                  .clk             ( clk                         ),
                  .rst_n           ( rst_n                       ),
                  .icache_is_private_i ( 1'b1                    ),
                  .test_en_i       ( test_en_i                   ),

                  // ---------------------------------------------------------------
                  // SHARED_ICACHE_INTERCONNECT Port Declarations -----------------------------------------
                  // ---------------------------------------------------------------
                  .fetch_req_i     (  instr_req_FB_to_IC[i]      ),
                  .fetch_grant_o   (  instr_gnt_FB_to_IC[i]      ),
                  .fetch_addr_i    (  instr_add_FB_to_IC[i]      ),
                  .fetch_ID_i      (  '0                         ),
                  .fetch_r_rdata_o (  instr_r_rdata_FB_to_IC[i]  ),
                  .fetch_r_valid_o (  instr_r_valid_FB_to_IC[i]  ),
                  .fetch_r_ID_o    (                             ),

                  // §§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§ //
                  // §§§§§§§§§§§§§§§§§§§    REFILL Request side  §§§§§§§§§§§§§§§§§§§§§§§ //
                  // §§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§§ //

                  .init_awid_o     (  init_awid_internal[i]     ),
                  .init_awaddr_o   (  init_awaddr_internal[i]   ),
                  .init_awlen_o    (  init_awlen_internal[i]    ),
                  .init_awsize_o   (  init_awsize_internal[i]   ),
                  .init_awburst_o  (  init_awburst_internal[i]  ),
                  .init_awlock_o   (  init_awlock_internal[i]   ),
                  .init_awcache_o  (  init_awcache_internal[i]  ),
                  .init_awprot_o   (  init_awprot_internal[i]   ),
                  .init_awregion_o (  init_awregion_internal[i] ),
                  .init_awuser_o   (  init_awuser_internal[i]   ),
                  .init_awqos_o    (  init_awqos_internal[i]    ),
                  .init_awvalid_o  (  init_awvalid_internal[i]  ),
                  .init_awready_i  (  init_awready_internal[i]  ),

                  .init_wdata_o    (  init_wdata_internal[i]    ),
                  .init_wstrb_o    (  init_wstrb_internal[i]    ),
                  .init_wlast_o    (  init_wlast_internal[i]    ),
                  .init_wuser_o    (  init_wuser_internal[i]    ),
                  .init_wvalid_o   (  init_wvalid_internal[i]   ),
                  .init_wready_i   (  init_wready_internal[i]   ),



                  .init_bid_i      (  init_bid_internal[i]      ),
                  .init_bresp_i    (  init_bresp_internal[i]    ),
                  .init_buser_i    (  init_buser_internal[i]    ),
                  .init_bvalid_i   (  init_bvalid_internal[i]   ),
                  .init_bready_o   (  init_bready_internal[i]   ),


                  .init_arid_o     (  init_arid_internal[i]     ),
                  .init_araddr_o   (  init_araddr_internal[i]   ),
                  .init_arlen_o    (  init_arlen_internal[i]    ),
                  .init_arsize_o   (  init_arsize_internal[i]   ),
                  .init_arburst_o  (  init_arburst_internal[i]  ),
                  .init_arlock_o   (  init_arlock_internal[i]   ),
                  .init_arcache_o  (  init_arcache_internal[i]  ),
                  .init_arprot_o   (  init_arprot_internal[i]   ),
                  .init_arregion_o (  init_arregion_internal[i] ),
                  .init_aruser_o   (  init_aruser_internal[i]   ),
                  .init_arqos_o    (  init_arqos_internal[i]    ),
                  .init_arvalid_o  (  init_arvalid_internal[i]  ),
                  .init_arready_i  (  init_arready_internal[i]  ),

                  .init_rid_i     (  init_rid_internal[i]       ),
                  .init_rdata_i   (  init_rdata_internal[i]     ),
                  .init_rresp_i   (  init_rresp_internal[i]     ),
                  .init_rlast_i   (  init_rlast_internal[i]     ),
                  .init_ruser_i   (  init_ruser_internal[i]     ),
                  .init_rvalid_i  (  init_rvalid_internal[i]    ),
                  .init_rready_o  (  init_rready_internal[i]    ),

                  // Control ports
                  .ctrl_req_enable_icache_i      ( IC_ctrl_unit_slave_if[i].ctrl_req_enable    ),
                  .ctrl_ack_enable_icache_o      ( IC_ctrl_unit_slave_if[i].ctrl_ack_enable    ),
                  .ctrl_req_disable_icache_i     ( IC_ctrl_unit_slave_if[i].ctrl_req_disable   ),
                  .ctrl_ack_disable_icache_o     ( IC_ctrl_unit_slave_if[i].ctrl_ack_disable   ),
                  .ctrl_pending_trans_icache_o   ( IC_ctrl_unit_slave_if[i].ctrl_pending_trans )
      `ifdef FEATURE_ICACHE_STAT
                  ,
                  .ctrl_hit_count_icache_o       ( IC_ctrl_unit_slave_if[i].ctrl_hit_count     ),
                  .ctrl_trans_count_icache_o     ( IC_ctrl_unit_slave_if[i].ctrl_trans_count   ),
                  .ctrl_clear_regs_icache_i      ( IC_ctrl_unit_slave_if[i].ctrl_clear_regs    ),
                  .ctrl_enable_regs_icache_i     ( IC_ctrl_unit_slave_if[i].ctrl_enable_regs   )
      `endif
                );

            end

  end
endgenerate

// fconti: workaround because Vivado synthesizes the '1 SystemVerilog construct
//         as LSB to 1 and other bits to 0, instead of all bits to 1

  logic [NB_REFILL_PORT-1:0][32-1:0]             axi_instr_bus_init_START_ADDR;
  logic [NB_REFILL_PORT-1:0][32-1:0]             axi_instr_bus_init_END_ADDR;
  logic [NB_REFILL_PORT-1:0]                     axi_instr_bus_init_valid_rule;
  `ifdef PRIVATE_ICACHE
  logic [NB_CORES-1:0][NB_REFILL_PORT-1:0] axi_instr_bus_init_connectivity_map; //FIXME
  `else
  logic [NB_CACHE_BANKS-1:0][NB_REFILL_PORT-1:0]       axi_instr_bus_init_connectivity_map; //FIXME
  `endif

  assign axi_instr_bus_init_START_ADDR = {NB_REFILL_PORT{32'h0}};
  assign axi_instr_bus_init_END_ADDR   = {NB_REFILL_PORT{32'hffffffff}};
  assign axi_instr_bus_init_valid_rule = {NB_REFILL_PORT{1'b1}};
  `ifdef PRIVATE_ICACHE
  assign axi_instr_bus_init_connectivity_map = {NB_CORES*NB_REFILL_PORT{1'b1}};//FIXME
  `else
  assign axi_instr_bus_init_connectivity_map = {NB_CACHE_BANKS*NB_REFILL_PORT{1'b1}};//FIXME
  `endif




/////////////////////////////////////////////////////////////////
//  █████╗ ██╗  ██╗██╗    ███╗   ██╗ ██████╗ ██████╗ ███████╗  //
// ██╔══██╗╚██╗██╔╝██║    ████╗  ██║██╔═══██╗██╔══██╗██╔════╝  //
// ███████║ ╚███╔╝ ██║    ██╔██╗ ██║██║   ██║██║  ██║█████╗    //
// ██╔══██║ ██╔██╗ ██║    ██║╚██╗██║██║   ██║██║  ██║██╔══╝    //
// ██║  ██║██╔╝ ██╗██║    ██║ ╚████║╚██████╔╝██████╔╝███████╗  //
// ╚═╝  ╚═╝╚═╝  ╚═╝╚═╝    ╚═╝  ╚═══╝ ╚═════╝ ╚═════╝ ╚══════╝  //
/////////////////////////////////////////////////////////////////
axi_node
#(

    .AXI_ADDRESS_W      ( AXI_ADDR       ),
    .AXI_DATA_W         ( AXI_DATA       ),
    .AXI_NUMBYTES       ( AXI_DATA/8     ),

    .AXI_USER_W         ( AXI_USER       ),
    .AXI_ID_IN          ( AXI_ID_INT     ),
    .AXI_ID_OUT         ( AXI_ID_OUT     ),

    .N_MASTER_PORT      ( NB_REFILL_PORT ),
    .N_SLAVE_PORT       ( NB_CACHE_BANKS ),


    .FIFO_DEPTH_DW      ( 2              ),
    .N_REGION           ( 1              )
)
AXI_INTRUCTION_BUS
(
  .clk                  (  clk                    ),
  .rst_n                (  rst_n                  ),
  .test_en_i            (  test_en_i              ),

  // ---------------------------------------------------------------
  // AXI TARG Port Declarations -----------------------------------------
  // ---------------------------------------------------------------
  .slave_awid_i          ( init_awid_internal      ),
  .slave_awaddr_i        ( init_awaddr_internal    ),
  .slave_awlen_i         ( init_awlen_internal     ),
  .slave_awsize_i        ( init_awsize_internal    ),
  .slave_awburst_i       ( init_awburst_internal   ),
  .slave_awlock_i        ( init_awlock_internal    ),
  .slave_awcache_i       ( init_awcache_internal   ),
  .slave_awprot_i        ( init_awprot_internal    ),
  .slave_awregion_i      ( init_awregion_internal  ),
  .slave_awuser_i        ( init_awuser_internal    ),
  .slave_awqos_i         ( init_awqos_internal     ),
  .slave_awvalid_i       ( init_awvalid_internal   ),
  .slave_awready_o       ( init_awready_internal   ),

  .slave_wdata_i         ( init_wdata_internal     ),
  .slave_wstrb_i         ( init_wstrb_internal     ),
  .slave_wlast_i         ( init_wlast_internal     ),
  .slave_wuser_i         ( init_wuser_internal     ),
  .slave_wvalid_i        ( init_wvalid_internal    ),
  .slave_wready_o        ( init_wready_internal    ),


  .slave_bid_o           ( init_bid_internal       ),
  .slave_bresp_o         ( init_bresp_internal     ),
  .slave_bvalid_o        ( init_bvalid_internal    ),
  .slave_buser_o         ( init_buser_internal     ),
  .slave_bready_i        ( init_bready_internal    ),


  .slave_arid_i          ( init_arid_internal      ),
  .slave_araddr_i        ( init_araddr_internal    ),
  .slave_arlen_i         ( init_arlen_internal     ),
  .slave_arsize_i        ( init_arsize_internal    ),
  .slave_arburst_i       ( init_arburst_internal   ),
  .slave_arlock_i        ( init_arlock_internal    ),
  .slave_arcache_i       ( init_arcache_internal   ),
  .slave_arprot_i        ( init_arprot_internal    ),
  .slave_arregion_i      ( init_arregion_internal  ),
  .slave_aruser_i        ( init_aruser_internal    ),
  .slave_arqos_i         ( init_arqos_internal     ),
  .slave_arvalid_i       ( init_arvalid_internal   ),
  .slave_arready_o       ( init_arready_internal   ),
  // -----------------------------------------------

  .slave_rid_o           ( init_rid_internal       ),
  .slave_rdata_o         ( init_rdata_internal     ),
  .slave_rresp_o         ( init_rresp_internal     ),
  .slave_rlast_o         ( init_rlast_internal     ),
  .slave_ruser_o         ( init_ruser_internal     ),
  .slave_rvalid_o        ( init_rvalid_internal    ),
  .slave_rready_i        ( init_rready_internal    ),
  // -----------------------------------------------

  // -----------------------------------------------
  // AXI INIT Port Declarations --------------------
  // -----------------------------------------------
  .master_awid_o          ( init_awid_o[AXI_ID_OUT-1:0] ),
  .master_awaddr_o        ( init_awaddr_o               ),
  .master_awlen_o         ( init_awlen_o                ),
  .master_awsize_o        ( init_awsize_o               ),
  .master_awburst_o       ( init_awburst_o              ),
  .master_awlock_o        ( init_awlock_o               ),
  .master_awcache_o       ( init_awcache_o              ),
  .master_awprot_o        ( init_awprot_o               ),
  .master_awregion_o      ( init_awregion_o             ),
  .master_awuser_o        ( init_awuser_o               ),
  .master_awqos_o         ( init_awqos_o                ),
  .master_awvalid_o       ( init_awvalid_o              ),
  .master_awready_i       ( init_awready_i              ),

  .master_wdata_o         ( init_wdata_o                ),
  .master_wstrb_o         ( init_wstrb_o                ),
  .master_wlast_o         ( init_wlast_o                ),
  .master_wuser_o         ( init_wuser_o                ),
  .master_wvalid_o        ( init_wvalid_o               ),
  .master_wready_i        ( init_wready_i               ),

  .master_bid_i           ( init_bid_i[AXI_ID_OUT-1:0]  ),
  .master_bresp_i         ( init_bresp_i                ),
  .master_buser_i         ( init_buser_i                ),
  .master_bvalid_i        ( init_bvalid_i               ),
  .master_bready_o        ( init_bready_o               ),

  .master_arid_o          ( init_arid_o[AXI_ID_OUT-1:0] ),
  .master_araddr_o        ( init_araddr_o               ),
  .master_arlen_o         ( init_arlen_o                ),
  .master_arsize_o        ( init_arsize_o               ),
  .master_arburst_o       ( init_arburst_o              ),
  .master_arlock_o        ( init_arlock_o               ),
  .master_arcache_o       ( init_arcache_o              ),
  .master_arprot_o        ( init_arprot_o               ),
  .master_arregion_o      ( init_arregion_o             ),
  .master_aruser_o        ( init_aruser_o               ),
  .master_arqos_o         ( init_arqos_o                ),
  .master_arvalid_o       ( init_arvalid_o              ),
  .master_arready_i       ( init_arready_i              ),

  .master_rid_i           ( init_rid_i[AXI_ID_OUT-1:0]  ),
  .master_rdata_i         ( init_rdata_i                ),
  .master_rresp_i         ( init_rresp_i                ),
  .master_rlast_i         ( init_rlast_i                ),
  .master_ruser_i         ( init_ruser_i                ),
  .master_rvalid_i        ( init_rvalid_i               ),
  .master_rready_o        ( init_rready_o               ),

  //Initial Memory map
  // fconti: workaround because Vivado synthesizes the '1 SystemVerilog construct
  //         as LSB to 1 and other bits to 0, instead of all bits to 1

  .cfg_START_ADDR_i       (axi_instr_bus_init_START_ADDR      ),
  .cfg_END_ADDR_i         (axi_instr_bus_init_END_ADDR        ),
  .cfg_valid_rule_i       (axi_instr_bus_init_valid_rule      ),
  .cfg_connectivity_map_i (axi_instr_bus_init_connectivity_map)


);

assign     init_awid_o[AXI_ID-1:AXI_ID_OUT] = '0;
assign     init_arid_o[AXI_ID-1:AXI_ID_OUT] = '0;



//------------------------------------------------------------------------------------------//
// ██████╗  █████╗ ██████╗  █████╗ ███╗   ███╗     ██████╗██╗  ██╗███████╗ ██████╗██╗  ██╗  //
// ██╔══██╗██╔══██╗██╔══██╗██╔══██╗████╗ ████║    ██╔════╝██║  ██║██╔════╝██╔════╝██║ ██╔╝  //
// ██████╔╝███████║██████╔╝███████║██╔████╔██║    ██║     ███████║█████╗  ██║     █████╔╝   //
// ██╔═══╝ ██╔══██║██╔══██╗██╔══██║██║╚██╔╝██║    ██║     ██╔══██║██╔══╝  ██║     ██╔═██╗   //
// ██║     ██║  ██║██║  ██║██║  ██║██║ ╚═╝ ██║    ╚██████╗██║  ██║███████╗╚██████╗██║  ██╗  //
// ╚═╝     ╚═╝  ╚═╝╚═╝  ╚═╝╚═╝  ╚═╝╚═╝     ╚═╝     ╚═════╝╚═╝  ╚═╝╚══════╝ ╚═════╝╚═╝  ╚═╝  //
//------------------------------------------------------------------------------------------//

//synopsys translate_off
initial
begin

     if(NB_REFILL_PORT != 1)
       $fatal(2,"NB_REFILL_PORT OUT OF ALLOWED RANGES");

     if( 2**`log2(CACHE_SIZE-1) != CACHE_SIZE)
        $fatal(2,"Icahe capacity not power of 2");

     if( (ICACHE_DATA_WIDTH < 32 ) || (2**`log2(ICACHE_DATA_WIDTH-1) != ICACHE_DATA_WIDTH) )
        $fatal(2,"ICACHE_DATA_WIDTH OUT OF ALLOWED RANGES");

     // CHECK POWER OF 2 parameters
     if( (2**`log2(CACHE_LINE-1) != CACHE_LINE) )
     begin : _CHECK_CACHE_LINE_POWER_2
         $fatal(2,"CACHE LINE  NOT POWER OF TWO");
     end

      // CHECK POWER OF 2 parameters
     if( (SET_ASSOCIATIVE < 1) || (2**`log2(SET_ASSOCIATIVE-1) != SET_ASSOCIATIVE) )
     begin : _CHECK_SET_ASSOCIATIVE_
         $fatal(2,"SET_ASSOCIATIVE OUT OF ALLOWED RANGES");
     end


     if(`log2(NB_CORES-1)+`log2(NB_CACHE_BANKS-1) > AXI_ID+1 )
     begin : _CHECK_ID_OVERFLOW_
         $fatal(2,"AXI ID OVERFLOW");
     end

     if( (NB_CORES < 1)  || (NB_CORES > 32) || (2**`log2(NB_CORES-1) != NB_CORES) )
     begin : _CHECK_NB_CORES_
         $fatal(2,"NUMBER OF CORES NOT COMPATIBLE");
     end

     if( (NB_CACHE_BANKS < 1)  || (NB_CACHE_BANKS > 32) || (2**`log2(NB_CACHE_BANKS-1) != NB_CACHE_BANKS) )
     begin : _CHECK_NB_CACHE_BANKS_
         $fatal(2,"NUMBER OF CACHE_BANKS NOT COMPATIBLE");
     end

     if(CACHE_LINE*ICACHE_DATA_WIDTH < 64)
     begin : _CHECK_CACHE_LINE_WIDTH_
         $fatal(2,"CACHE LINE SIZE (%d bits) MUST BE >= 64bits", CACHE_LINE*ICACHE_DATA_WIDTH);
     end

     if((L0_SIZE != ICACHE_DATA_WIDTH) && (L0_BUFFER_FEATURE == "ENABLED"))
     begin : _CHECK_L0_SIZE
         $fatal(2,"L0_BUFFER SIZE and ICACHE_DATA_WIDTH MISMATCH", L0_SIZE, ICACHE_DATA_WIDTH);
     end

     if( ~((DIRECT_MAPPED_FEATURE == "ENABLED") || (DIRECT_MAPPED_FEATURE == "DISABLED"))  )
     begin : _CHECK_DIRECT_MAPPED_FEATURE_VALUE
         $fatal(2,"DIRECT_MAPPED_FEATURE can be DISABLED or ENABLED only. Passed %s. Please Correct it!", DIRECT_MAPPED_FEATURE );
     end

     if( (DIRECT_MAPPED_FEATURE == "ENABLED") &&  ( SET_ASSOCIATIVE > 1) )
     begin : _CHECK_DIRECT_MAPPED_VS_SET_ASSOCIATIVE_
         $fatal(2,"CACHE CONFIGURED AS DIRECT MAPPED (%s), WHILE NUMBER OF WAY is > 1 (%d)!", DIRECT_MAPPED_FEATURE, SET_ASSOCIATIVE );
     end

     if((ICACHE_DATA_WIDTH > 32)  && (L0_BUFFER_FEATURE == "DISABLED") && (ICACHE_DATA_WIDTH != INSTR_RDATA_WIDTH))
     begin : _CHECK_L0_ENABLED_
        $fatal(2,"ICACHE_DATA_WIDTH is (%d) and not equal to INSTR_RDATA_WIDTH (%d) and thus requires an enabled L0_BUFFER (%s)", ICACHE_DATA_WIDTH, INSTR_RDATA_WIDTH, L0_BUFFER_FEATURE );
     end

     if((L0_BUFFER_FEATURE == "ENABLED") && (INSTR_RDATA_WIDTH != 32))
     begin : _CHECK_L0_ENABLED_INSTR_RDATA
        $fatal(2,"INSTR_RDATA_WIDTH is (%d) and L0_BUFFER is enabled (%s), INSTR_RDATA_WIDTH needs to be 32", L0_BUFFER_FEATURE, INSTR_RDATA_WIDTH );
     end


    if(SHARED_ICACHE == "DISABLED")
    begin : CHECK_PRIVATE_CACHES
        if(NB_CORES != NB_CACHE_BANKS)
          $fatal(2,"Private cache Error: istantiated %d Cache banks with %d CORES", NB_CACHE_BANKS, NB_CORES);

        if((CACHE_SIZE*8)/(ICACHE_DATA_WIDTH*CACHE_LINE) == 1)
          $error("TAGRAM too SMALL (2 rows only)", NB_CACHE_BANKS, NB_CORES);
    end
    else
    begin : CHECK_SHARED_CACHES
        if((CACHE_SIZE*8)/(NB_CACHE_BANKS*ICACHE_DATA_WIDTH*CACHE_LINE) == 1)
          $error("TAGRAM too SMALL (2 row only)", NB_CACHE_BANKS, NB_CORES);
    end

end
//synopsys translate_on
endmodule
