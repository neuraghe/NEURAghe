// SOC BUS PARAMETRES
`include "ulpsoc_defines.sv"

`define NB_SLAVE  2
`define NB_MASTER 6


`define NB_REGION 1


    // MASTER PORT TO CORE MEM
    `define MASTER_0_START_ADDR 32'h1000_0000
    `define MASTER_0_END_ADDR   32'h1000_7FFF
    
    // MASTER PORT TO L3 via RAB
    `define MASTER_1_START_ADDR 32'h8000_0000
    `define MASTER_1_END_ADDR   32'hFFFF_FFFF

    // MASTER PORT TO L2(64MB)
    `define MASTER_2_START_ADDR 32'h1C00_0000
    `define MASTER_2_END_ADDR   32'h1FFF_FFFF

    // MASTER PORT TO STDOUT(64KB)
    `define MASTER_3_START_ADDR 32'h1A11_0000
    `define MASTER_3_END_ADDR   32'h1A11_FFFF    

    // MASTER PORT TO PERIPHERAL INTERCONNECT
    `define MASTER_4_START_ADDR 32'h1020_0000
    `define MASTER_4_END_ADDR   32'h102F_FFFF

    // MASTER PORT TO WEIGHTS DMA
    `define MASTER_5_START_ADDR 32'h1030_0000
    `define MASTER_5_END_ADDR   32'h103F_FFFF
