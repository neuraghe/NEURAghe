// CLUSTER BUS PARAMETRES

`define NB_SLAVE  4
`define NB_MASTER 4

`define NB_REGION 1

// MSTER PORT TO TCDM
`define MASTER_0_START_ADDR 32'h1000_0000
`define MASTER_0_END_ADDR   32'h101F_FFFF

// MASTER PORT TO PERIPHERAL INTERCONNECT
`define MASTER_1_START_ADDR 32'h1020_0000
`define MASTER_1_END_ADDR   32'h102F_FFFF

// MASTER PORT TO SOC (SOC PERIPHERALS + L2)
`define MASTER_2_START_ADDR 32'h1A00_0000
`define MASTER_2_END_ADDR   32'hFFFF_FFFF

// MASTER PORT TO WEIGHTS DMA
`define MASTER_3_START_ADDR 32'h1030_0000
`define MASTER_3_END_ADDR   32'h103F_FFFF
