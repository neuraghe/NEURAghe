`timescale 1ns/1ps

`celldefine
module AD42M2RA( CO, ICO, S, A, B, C, D, ICI);
input A, B, C, D, ICI;
output CO, ICO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AD42M2RA$func AD42M2RA_inst(.A(A),.B(B),.C(C),.CO(CO),.D(D),.ICI(ICI),.ICO(ICO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AD42M2RA$func AD42M2RA_inst(.A(A),.B(B),.C(C),.CO(CO),.D(D),.ICI(ICI),.ICO(ICO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

        ifnone
	// arc posedge A --> (CO:A)
	 (posedge A => (CO:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (CO:A)
	 (negedge A => (CO:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

        ifnone
	// arc posedge B --> (CO:B)
	 (posedge B => (CO:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (CO:B)
	 (negedge B => (CO:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

        ifnone
	// arc posedge C --> (CO:C)
	 (posedge C => (CO:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (CO:C)
	 (negedge C => (CO:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	ifnone
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	ifnone
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	ifnone
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	ifnone
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	ifnone
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

        ifnone
	// arc posedge C --> (S:C)
	 (posedge C => (S:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (S:C)
	 (negedge C => (S:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

        ifnone
	// arc posedge D --> (S:D)
	 (posedge D => (S:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (S:D)
	 (negedge D => (S:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

        ifnone
	// arc posedge ICI --> (S:ICI)
	 (posedge ICI => (S:ICI)) = (1.0,1.0);

        ifnone
	// arc negedge ICI --> (S:ICI)
	 (negedge ICI => (S:ICI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AD42M4RA( CO, ICO, S, A, B, C, D, ICI);
input A, B, C, D, ICI;
output CO, ICO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AD42M4RA$func AD42M4RA_inst(.A(A),.B(B),.C(C),.CO(CO),.D(D),.ICI(ICI),.ICO(ICO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AD42M4RA$func AD42M4RA_inst(.A(A),.B(B),.C(C),.CO(CO),.D(D),.ICI(ICI),.ICO(ICO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

        ifnone
	// arc posedge A --> (CO:A)
	 (posedge A => (CO:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (CO:A)
	 (negedge A => (CO:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

        ifnone
	// arc posedge B --> (CO:B)
	 (posedge B => (CO:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (CO:B)
	 (negedge B => (CO:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

        ifnone
	// arc posedge C --> (CO:C)
	 (posedge C => (CO:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (CO:C)
	 (negedge C => (CO:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> CO
	 (C => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	ifnone
	// arc D --> CO
	 (D => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	ifnone
	// arc ICI --> CO
	 (ICI => CO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	ifnone
	// arc A --> ICO
	 (A => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	ifnone
	// arc B --> ICO
	 (B => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	ifnone
	// arc C --> ICO
	 (C => ICO) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

        ifnone
	// arc posedge C --> (S:C)
	 (posedge C => (S:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (S:C)
	 (negedge C => (S:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1)
	// arc C --> S
	 (C => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

        ifnone
	// arc posedge D --> (S:D)
	 (posedge D => (S:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (S:D)
	 (negedge D => (S:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1)
	// arc D --> S
	 (D => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

        ifnone
	// arc posedge ICI --> (S:ICI)
	 (posedge ICI => (S:ICI)) = (1.0,1.0);

        ifnone
	// arc negedge ICI --> (S:ICI)
	 (negedge ICI => (S:ICI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1)
	// arc ICI --> S
	 (ICI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADCSCM2R( CO0, CO1, A, B, NCI0, NCI1);
input A, B, NCI0, NCI1;
output CO0, CO1;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADCSCM2R$func ADCSCM2R_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.NCI0(NCI0),.NCI1(NCI1));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADCSCM2R$func ADCSCM2R_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.NCI0(NCI0),.NCI1(NCI1));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	ifnone
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	ifnone
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	ifnone
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	ifnone
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	ifnone
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	ifnone
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADCSCM4R( CO0, CO1, A, B, NCI0, NCI1);
input A, B, NCI0, NCI1;
output CO0, CO1;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADCSCM4R$func ADCSCM4R_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.NCI0(NCI0),.NCI1(NCI1));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADCSCM4R$func ADCSCM4R_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.NCI0(NCI0),.NCI1(NCI1));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	ifnone
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	ifnone
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	ifnone
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	ifnone
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	ifnone
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	ifnone
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADCSIOM2R( CO0B, CO1B, A, B);
input A, B;
output CO0B, CO1B;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADCSIOM2R$func ADCSIOM2R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADCSIOM2R$func ADCSIOM2R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADCSIOM4R( CO0B, CO1B, A, B);
input A, B;
output CO0B, CO1B;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADCSIOM4R$func ADCSIOM4R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADCSIOM4R$func ADCSIOM4R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADCSOM2R( CO0B, CO1B, A, B, CI0, CI1);
input A, B, CI0, CI1;
output CO0B, CO1B;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADCSOM2R$func ADCSOM2R_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADCSOM2R$func ADCSOM2R_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	ifnone
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	ifnone
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	ifnone
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	ifnone
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	ifnone
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	ifnone
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADCSOM4R( CO0B, CO1B, A, B, CI0, CI1);
input A, B, CI0, CI1;
output CO0B, CO1B;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADCSOM4R$func ADCSOM4R_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADCSOM4R$func ADCSOM4R_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	ifnone
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	ifnone
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	ifnone
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	ifnone
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	ifnone
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	ifnone
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCGCM2RA( CO, A, B, NCI);
input A, B, NCI;
output CO;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCGCM2RA$func ADFCGCM2RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCGCM2RA$func ADFCGCM2RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && NCI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	ifnone
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCGCM4RA( CO, A, B, NCI);
input A, B, NCI;
output CO;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCGCM4RA$func ADFCGCM4RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCGCM4RA$func ADFCGCM4RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && NCI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	ifnone
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCGOM2RA( COB, A, B, CI);
input A, B, CI;
output COB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCGOM2RA$func ADFCGOM2RA_inst(.A(A),.B(B),.CI(CI),.COB(COB));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCGOM2RA$func ADFCGOM2RA_inst(.A(A),.B(B),.CI(CI),.COB(COB));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	ifnone
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	ifnone
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	ifnone
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCGOM4RA( COB, A, B, CI);
input A, B, CI;
output COB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCGOM4RA$func ADFCGOM4RA_inst(.A(A),.B(B),.CI(CI),.COB(COB));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCGOM4RA$func ADFCGOM4RA_inst(.A(A),.B(B),.CI(CI),.COB(COB));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	ifnone
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	ifnone
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	ifnone
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCM2RA( CO, S, A, B, NCI);
input A, B, NCI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCM2RA$func ADFCM2RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCM2RA$func ADFCM2RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && NCI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	ifnone
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(B===1'b0 && NCI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

        ifnone
	// arc posedge NCI --> (S:NCI)
	 (posedge NCI => (S:NCI)) = (1.0,1.0);

        ifnone
	// arc negedge NCI --> (S:NCI)
	 (negedge NCI => (S:NCI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCM4RA( CO, S, A, B, NCI);
input A, B, NCI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCM4RA$func ADFCM4RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCM4RA$func ADFCM4RA_inst(.A(A),.B(B),.CO(CO),.NCI(NCI),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && NCI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	ifnone
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(B===1'b0 && NCI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && NCI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && NCI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && NCI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

        ifnone
	// arc posedge NCI --> (S:NCI)
	 (posedge NCI => (S:NCI)) = (1.0,1.0);

        ifnone
	// arc negedge NCI --> (S:NCI)
	 (negedge NCI => (S:NCI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc NCI --> S
	 (NCI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCSCM2RA( CO0, CO1, S, A, B, CS, NCI0, NCI1);
input A, B, CS, NCI0, NCI1;
output CO0, CO1, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCSCM2RA$func ADFCSCM2RA_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.CS(CS),.NCI0(NCI0),.NCI1(NCI1),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCSCM2RA$func ADFCSCM2RA_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.CS(CS),.NCI0(NCI0),.NCI1(NCI1),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	ifnone
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	ifnone
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	ifnone
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	ifnone
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	ifnone
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	ifnone
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

        ifnone
	// arc posedge NCI0 --> (S:NCI0)
	 (posedge NCI0 => (S:NCI0)) = (1.0,1.0);

        ifnone
	// arc negedge NCI0 --> (S:NCI0)
	 (negedge NCI0 => (S:NCI0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

        ifnone
	// arc posedge NCI1 --> (S:NCI1)
	 (posedge NCI1 => (S:NCI1)) = (1.0,1.0);

        ifnone
	// arc negedge NCI1 --> (S:NCI1)
	 (negedge NCI1 => (S:NCI1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCSCM4RA( CO0, CO1, S, A, B, CS, NCI0, NCI1);
input A, B, CS, NCI0, NCI1;
output CO0, CO1, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCSCM4RA$func ADFCSCM4RA_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.CS(CS),.NCI0(NCI0),.NCI1(NCI1),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCSCM4RA$func ADFCSCM4RA_inst(.A(A),.B(B),.CO0(CO0),.CO1(CO1),.CS(CS),.NCI0(NCI0),.NCI1(NCI1),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	ifnone
	// arc A --> CO0
	 (A => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	ifnone
	// arc B --> CO0
	 (B => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b0)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b1)
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	ifnone
	// arc NCI0 --> CO0
	 (NCI0 => CO0) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	ifnone
	// arc A --> CO1
	 (A => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	ifnone
	// arc B --> CO1
	 (B => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	ifnone
	// arc NCI1 --> CO1
	 (NCI1 => CO1) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

        ifnone
	// arc posedge NCI0 --> (S:NCI0)
	 (posedge NCI0 => (S:NCI0)) = (1.0,1.0);

        ifnone
	// arc negedge NCI0 --> (S:NCI0)
	 (negedge NCI0 => (S:NCI0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b0)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI1===1'b1)
	// arc NCI0 --> S
	 (NCI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

        ifnone
	// arc posedge NCI1 --> (S:NCI1)
	 (posedge NCI1 => (S:NCI1)) = (1.0,1.0);

        ifnone
	// arc negedge NCI1 --> (S:NCI1)
	 (negedge NCI1 => (S:NCI1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b0)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && NCI0===1'b1)
	// arc NCI1 --> S
	 (NCI1 => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCSIOM2R( CO0B, CO1B, S, A, B, CS);
input A, B, CS;
output CO0B, CO1B, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCSIOM2R$func ADFCSIOM2R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCSIOM2R$func ADFCSIOM2R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	ifnone
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	ifnone
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	ifnone
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	ifnone
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCSIOM4R( CO0B, CO1B, S, A, B, CS);
input A, B, CS;
output CO0B, CO1B, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCSIOM4R$func ADFCSIOM4R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCSIOM4R$func ADFCSIOM4R_inst(.A(A),.B(B),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	ifnone
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	ifnone
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	ifnone
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	ifnone
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(B===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCSOM2RA( CO0B, CO1B, S, A, B, CI0, CI1, CS);
input A, B, CI0, CI1, CS;
output CO0B, CO1B, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCSOM2RA$func ADFCSOM2RA_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCSOM2RA$func ADFCSOM2RA_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	ifnone
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	ifnone
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	ifnone
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	ifnone
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	ifnone
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	ifnone
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

        ifnone
	// arc posedge CI0 --> (S:CI0)
	 (posedge CI0 => (S:CI0)) = (1.0,1.0);

        ifnone
	// arc negedge CI0 --> (S:CI0)
	 (negedge CI0 => (S:CI0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

        ifnone
	// arc posedge CI1 --> (S:CI1)
	 (posedge CI1 => (S:CI1)) = (1.0,1.0);

        ifnone
	// arc negedge CI1 --> (S:CI1)
	 (negedge CI1 => (S:CI1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFCSOM4RA( CO0B, CO1B, S, A, B, CI0, CI1, CS);
input A, B, CI0, CI1, CS;
output CO0B, CO1B, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFCSOM4RA$func ADFCSOM4RA_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFCSOM4RA$func ADFCSOM4RA_inst(.A(A),.B(B),.CI0(CI0),.CI1(CI1),.CO0B(CO0B),.CO1B(CO1B),.CS(CS),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	ifnone
	// arc A --> CO0B
	 (A => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	ifnone
	// arc B --> CO0B
	 (B => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	ifnone
	// arc CI0 --> CO0B
	 (CI0 => CO0B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	ifnone
	// arc A --> CO1B
	 (A => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	ifnone
	// arc B --> CO1B
	 (B => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b0)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1)
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	ifnone
	// arc CI1 --> CO1B
	 (CI1 => CO1B) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

        ifnone
	// arc posedge CI0 --> (S:CI0)
	 (posedge CI0 => (S:CI0)) = (1.0,1.0);

        ifnone
	// arc negedge CI0 --> (S:CI0)
	 (negedge CI0 => (S:CI0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI1===1'b0)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI1===1'b1)
	// arc CI0 --> S
	 (CI0 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

        ifnone
	// arc posedge CI1 --> (S:CI1)
	 (posedge CI1 => (S:CI1)) = (1.0,1.0);

        ifnone
	// arc negedge CI1 --> (S:CI1)
	 (negedge CI1 => (S:CI1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b0)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b1)
	// arc CI1 --> S
	 (CI1 => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
	// arc CS --> S
	 (CS => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFM0RA( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFM0RA$func ADFM0RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFM0RA$func ADFM0RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFM1RA( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFM1RA$func ADFM1RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFM1RA$func ADFM1RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFM2RA( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFM2RA$func ADFM2RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFM2RA$func ADFM2RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFM4RA( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFM4RA$func ADFM4RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFM4RA$func ADFM4RA_inst(.A(A),.B(B),.CI(CI),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	ifnone
	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	ifnone
	// arc CI --> CO
	 (CI => CO) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFOM2RA( COB, S, A, B, CI);
input A, B, CI;
output COB, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFOM2RA$func ADFOM2RA_inst(.A(A),.B(B),.CI(CI),.COB(COB),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFOM2RA$func ADFOM2RA_inst(.A(A),.B(B),.CI(CI),.COB(COB),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	ifnone
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	ifnone
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	ifnone
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADFOM4RA( COB, S, A, B, CI);
input A, B, CI;
output COB, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADFOM4RA$func ADFOM4RA_inst(.A(A),.B(B),.CI(CI),.COB(COB),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADFOM4RA$func ADFOM4RA_inst(.A(A),.B(B),.CI(CI),.COB(COB),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && CI===1'b1)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	ifnone
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	ifnone
	// arc B --> COB
	 (B => COB) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	ifnone
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(B===1'b0 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(B===1'b0 && CI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(B===1'b1 && CI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(A===1'b0 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

        ifnone
	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

	if(A===1'b0 && CI===1'b0)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b1 && CI===1'b1)
	// arc B --> S
	 (B => S) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc CI --> S
	 (CI => S) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHCM2R( CO, S, A, NCI);
input A, NCI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHCM2R$func ADHCM2R_inst(.A(A),.CO(CO),.NCI(NCI),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHCM2R$func ADHCM2R_inst(.A(A),.CO(CO),.NCI(NCI),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge NCI --> (S:NCI)
	 (posedge NCI => (S:NCI)) = (1.0,1.0);

	// arc negedge NCI --> (S:NCI)
	 (negedge NCI => (S:NCI)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHCM4R( CO, S, A, NCI);
input A, NCI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHCM4R$func ADHCM4R_inst(.A(A),.CO(CO),.NCI(NCI),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHCM4R$func ADHCM4R_inst(.A(A),.CO(CO),.NCI(NCI),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge NCI --> (S:NCI)
	 (posedge NCI => (S:NCI)) = (1.0,1.0);

	// arc negedge NCI --> (S:NCI)
	 (negedge NCI => (S:NCI)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHCSCM2R( CO, S, A, CS, NCI);
input A, CS, NCI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHCSCM2R$func ADHCSCM2R_inst(.A(A),.CO(CO),.CS(CS),.NCI(NCI),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHCSCM2R$func ADHCSCM2R_inst(.A(A),.CO(CO),.CS(CS),.NCI(NCI),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(CS===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(CS===1'b0)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(CS===1'b1)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	ifnone
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(CS===1'b0 && NCI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CS===1'b0 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CS===1'b1 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc posedge NCI --> (S:NCI)
	 (posedge NCI => (S:NCI)) = (1.0,1.0);

        ifnone
	// arc negedge NCI --> (S:NCI)
	 (negedge NCI => (S:NCI)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHCSCM4R( CO, S, A, CS, NCI);
input A, CS, NCI;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHCSCM4R$func ADHCSCM4R_inst(.A(A),.CO(CO),.CS(CS),.NCI(NCI),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHCSCM4R$func ADHCSCM4R_inst(.A(A),.CO(CO),.CS(CS),.NCI(NCI),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(CS===1'b0)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	ifnone
	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	if(CS===1'b0)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	if(CS===1'b1)
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

	ifnone
	// arc NCI --> CO
	 (NCI => CO) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(CS===1'b0 && NCI===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CS===1'b0 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CS===1'b1 && NCI===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc posedge NCI --> (S:NCI)
	 (posedge NCI => (S:NCI)) = (1.0,1.0);

        ifnone
	// arc negedge NCI --> (S:NCI)
	 (negedge NCI => (S:NCI)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHCSOM2R( COB, S, A, CI, CS);
input A, CI, CS;
output COB, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHCSOM2R$func ADHCSOM2R_inst(.A(A),.CI(CI),.COB(COB),.CS(CS),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHCSOM2R$func ADHCSOM2R_inst(.A(A),.CI(CI),.COB(COB),.CS(CS),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(CS===1'b0)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	ifnone
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(CS===1'b0)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(CS===1'b1)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	ifnone
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(CI===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CI===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CI===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHCSOM4R( COB, S, A, CI, CS);
input A, CI, CS;
output COB, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHCSOM4R$func ADHCSOM4R_inst(.A(A),.CI(CI),.COB(COB),.CS(CS),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHCSOM4R$func ADHCSOM4R_inst(.A(A),.CI(CI),.COB(COB),.CS(CS),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(CS===1'b0)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(CS===1'b1)
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	ifnone
	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	if(CS===1'b0)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	if(CS===1'b1)
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	ifnone
	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

        ifnone
	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	if(CI===1'b0 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CI===1'b0 && CS===1'b1)
	// arc A --> S
	 (A => S) = (1.0,1.0);

	if(CI===1'b1 && CS===1'b0)
	// arc A --> S
	 (A => S) = (1.0,1.0);

        ifnone
	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

        ifnone
	// arc posedge CS --> (S:CS)
	 (posedge CS => (S:CS)) = (1.0,1.0);

        ifnone
	// arc negedge CS --> (S:CS)
	 (negedge CS => (S:CS)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHM1RA( CO, S, A, B);
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHM1RA$func ADHM1RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHM1RA$func ADHM1RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHM2RA( CO, S, A, B);
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHM2RA$func ADHM2RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHM2RA$func ADHM2RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHM4RA( CO, S, A, B);
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHM4RA$func ADHM4RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHM4RA$func ADHM4RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHM8RA( CO, S, A, B);
input A, B;
output CO, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHM8RA$func ADHM8RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHM8RA$func ADHM8RA_inst(.A(A),.B(B),.CO(CO),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> CO
	 (A => CO) = (1.0,1.0);

	// arc B --> CO
	 (B => CO) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge B --> (S:B)
	 (posedge B => (S:B)) = (1.0,1.0);

	// arc negedge B --> (S:B)
	 (negedge B => (S:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHOM2R( COB, S, A, CI);
input A, CI;
output COB, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHOM2R$func ADHOM2R_inst(.A(A),.CI(CI),.COB(COB),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHOM2R$func ADHOM2R_inst(.A(A),.CI(CI),.COB(COB),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ADHOM4R( COB, S, A, CI);
input A, CI;
output COB, S;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ADHOM4R$func ADHOM4R_inst(.A(A),.CI(CI),.COB(COB),.S(S));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ADHOM4R$func ADHOM4R_inst(.A(A),.CI(CI),.COB(COB),.S(S));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> COB
	 (A => COB) = (1.0,1.0);

	// arc CI --> COB
	 (CI => COB) = (1.0,1.0);

	// arc posedge A --> (S:A)
	 (posedge A => (S:A)) = (1.0,1.0);

	// arc negedge A --> (S:A)
	 (negedge A => (S:A)) = (1.0,1.0);

	// arc posedge CI --> (S:CI)
	 (posedge CI => (S:CI)) = (1.0,1.0);

	// arc negedge CI --> (S:CI)
	 (negedge CI => (S:CI)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M0R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M0R$func AN2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M0R$func AN2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M12RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M12RA$func AN2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M12RA$func AN2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M16RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M16RA$func AN2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M16RA$func AN2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M1R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M1R$func AN2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M1R$func AN2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M22RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M22RA$func AN2M22RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M22RA$func AN2M22RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M2R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M2R$func AN2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M2R$func AN2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M4R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M4R$func AN2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M4R$func AN2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M6R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M6R$func AN2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M6R$func AN2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN2M8R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN2M8R$func AN2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN2M8R$func AN2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M0R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M0R$func AN3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M0R$func AN3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M12RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M12RA$func AN3M12RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M12RA$func AN3M12RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M16RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M16RA$func AN3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M16RA$func AN3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M1R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M1R$func AN3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M1R$func AN3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M22RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M22RA$func AN3M22RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M22RA$func AN3M22RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M2R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M2R$func AN3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M2R$func AN3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M4R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M4R$func AN3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M4R$func AN3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M6R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M6R$func AN3M6R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M6R$func AN3M6R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN3M8R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN3M8R$func AN3M8R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN3M8R$func AN3M8R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M0R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M0R$func AN4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M0R$func AN4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M12RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M12RA$func AN4M12RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M12RA$func AN4M12RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M16RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M16RA$func AN4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M16RA$func AN4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M1R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M1R$func AN4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M1R$func AN4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M2R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M2R$func AN4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M2R$func AN4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M4RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M4RA$func AN4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M4RA$func AN4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M6R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M6R$func AN4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M6R$func AN4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AN4M8RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AN4M8RA$func AN4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AN4M8RA$func AN4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ANTR( A);
input A;

endmodule
`endcelldefine
`celldefine
module AO211M1RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO211M1RA$func AO211M1RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO211M1RA$func AO211M1RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO211M2RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO211M2RA$func AO211M2RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO211M2RA$func AO211M2RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO211M4RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO211M4RA$func AO211M4RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO211M4RA$func AO211M4RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO211M8RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO211M8RA$func AO211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO211M8RA$func AO211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M0RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M0RA$func AO21M0RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M0RA$func AO21M0RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M12RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M12RA$func AO21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M12RA$func AO21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M1RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M1RA$func AO21M1RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M1RA$func AO21M1RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M2RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M2RA$func AO21M2RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M2RA$func AO21M2RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M4RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M4RA$func AO21M4RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M4RA$func AO21M4RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M6RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M6RA$func AO21M6RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M6RA$func AO21M6RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO21M8RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO21M8RA$func AO21M8RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO21M8RA$func AO21M8RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO221M1RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO221M1RA$func AO221M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO221M1RA$func AO221M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO221M2RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO221M2RA$func AO221M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO221M2RA$func AO221M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO221M4RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO221M4RA$func AO221M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO221M4RA$func AO221M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO221M8RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO221M8RA$func AO221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO221M8RA$func AO221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO222M1RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO222M1RA$func AO222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO222M1RA$func AO222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO222M2RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO222M2RA$func AO222M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO222M2RA$func AO222M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO222M4RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO222M4RA$func AO222M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO222M4RA$func AO222M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO222M8RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO222M8RA$func AO222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO222M8RA$func AO222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B10M0R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B10M0R$func AO22B10M0R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B10M0R$func AO22B10M0R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B10M1R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B10M1R$func AO22B10M1R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B10M1R$func AO22B10M1R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B10M2R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B10M2R$func AO22B10M2R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B10M2R$func AO22B10M2R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B10M4R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B10M4R$func AO22B10M4R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B10M4R$func AO22B10M4R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B10M8RA( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B10M8RA$func AO22B10M8RA_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B10M8RA$func AO22B10M8RA_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B11M0R( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B11M0R$func AO22B11M0R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B11M0R$func AO22B11M0R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && NB2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B11M1R( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B11M1R$func AO22B11M1R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B11M1R$func AO22B11M1R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && NB2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B11M2R( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B11M2R$func AO22B11M2R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B11M2R$func AO22B11M2R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && NB2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B11M4R( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B11M4R$func AO22B11M4R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B11M4R$func AO22B11M4R_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && NB2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22B11M8RA( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22B11M8RA$func AO22B11M8RA_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22B11M8RA$func AO22B11M8RA_inst(.A1(A1),.B1(B1),.NA2(NA2),.NB2(NB2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && NB2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && NB2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

	ifnone
	// arc NB2 --> Z
	 (NB2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M0RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M0RA$func AO22M0RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M0RA$func AO22M0RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M12RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M12RA$func AO22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M12RA$func AO22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M1RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M1RA$func AO22M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M1RA$func AO22M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M2R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M2R$func AO22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M2R$func AO22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M4RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M4RA$func AO22M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M4RA$func AO22M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M6RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M6RA$func AO22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M6RA$func AO22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO22M8RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO22M8RA$func AO22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO22M8RA$func AO22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO31M1RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO31M1RA$func AO31M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO31M1RA$func AO31M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO31M2RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO31M2RA$func AO31M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO31M2RA$func AO31M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO31M4RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO31M4RA$func AO31M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO31M4RA$func AO31M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO31M8RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO31M8RA$func AO31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO31M8RA$func AO31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO32M1RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO32M1RA$func AO32M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO32M1RA$func AO32M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO32M2RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO32M2RA$func AO32M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO32M2RA$func AO32M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO32M4RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO32M4RA$func AO32M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO32M4RA$func AO32M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO32M8RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO32M8RA$func AO32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO32M8RA$func AO32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO33M1RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO33M1RA$func AO33M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO33M1RA$func AO33M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO33M2RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO33M2RA$func AO33M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO33M2RA$func AO33M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO33M4RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO33M4RA$func AO33M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO33M4RA$func AO33M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AO33M8RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AO33M8RA$func AO33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AO33M8RA$func AO33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI211M0R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI211M0R$func AOI211M0R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI211M0R$func AOI211M0R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI211M1R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI211M1R$func AOI211M1R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI211M1R$func AOI211M1R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI211M2R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI211M2R$func AOI211M2R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI211M2R$func AOI211M2R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI211M4R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI211M4R$func AOI211M4R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI211M4R$func AOI211M4R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI211M6RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI211M6RA$func AOI211M6RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI211M6RA$func AOI211M6RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI211M8RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI211M8RA$func AOI211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI211M8RA$func AOI211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M0R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M0R$func AOI21B01M0R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M0R$func AOI21B01M0R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M12RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M12RA$func AOI21B01M12RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M12RA$func AOI21B01M12RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M16RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M16RA$func AOI21B01M16RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M16RA$func AOI21B01M16RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M1R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M1R$func AOI21B01M1R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M1R$func AOI21B01M1R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M2R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M2R$func AOI21B01M2R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M2R$func AOI21B01M2R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M4R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M4R$func AOI21B01M4R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M4R$func AOI21B01M4R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M6RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M6RA$func AOI21B01M6RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M6RA$func AOI21B01M6RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B01M8RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B01M8RA$func AOI21B01M8RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B01M8RA$func AOI21B01M8RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M0R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M0R$func AOI21B10M0R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M0R$func AOI21B10M0R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M12RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M12RA$func AOI21B10M12RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M12RA$func AOI21B10M12RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M16RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M16RA$func AOI21B10M16RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M16RA$func AOI21B10M16RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M1R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M1R$func AOI21B10M1R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M1R$func AOI21B10M1R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M2R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M2R$func AOI21B10M2R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M2R$func AOI21B10M2R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M4R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M4R$func AOI21B10M4R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M4R$func AOI21B10M4R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M6RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M6RA$func AOI21B10M6RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M6RA$func AOI21B10M6RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B10M8RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B10M8RA$func AOI21B10M8RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B10M8RA$func AOI21B10M8RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B20M0R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B20M0R$func AOI21B20M0R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M0R$func AOI21B20M0R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B20M1R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B20M1R$func AOI21B20M1R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M1R$func AOI21B20M1R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B20M2R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B20M2R$func AOI21B20M2R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M2R$func AOI21B20M2R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B20M4R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B20M4R$func AOI21B20M4R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M4R$func AOI21B20M4R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21B20M8RA( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21B20M8RA$func AOI21B20M8RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21B20M8RA$func AOI21B20M8RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M0R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M0R$func AOI21M0R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M0R$func AOI21M0R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M12RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M12RA$func AOI21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M12RA$func AOI21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M16RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M16RA$func AOI21M16RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M16RA$func AOI21M16RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M1R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M1R$func AOI21M1R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M1R$func AOI21M1R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M2R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M2R$func AOI21M2R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M2R$func AOI21M2R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M3R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M3R$func AOI21M3R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M3R$func AOI21M3R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M4R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M4R$func AOI21M4R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M4R$func AOI21M4R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M6R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M6R$func AOI21M6R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M6R$func AOI21M6R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI21M8R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI21M8R$func AOI21M8R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI21M8R$func AOI21M8R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI221M0R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI221M0R$func AOI221M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI221M0R$func AOI221M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI221M1R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI221M1R$func AOI221M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI221M1R$func AOI221M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI221M2R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI221M2R$func AOI221M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI221M2R$func AOI221M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI221M4R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI221M4R$func AOI221M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI221M4R$func AOI221M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI221M6RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI221M6RA$func AOI221M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI221M6RA$func AOI221M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI221M8RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI221M8RA$func AOI221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI221M8RA$func AOI221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI222M0RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI222M0RA$func AOI222M0RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI222M0RA$func AOI222M0RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI222M1RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI222M1RA$func AOI222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI222M1RA$func AOI222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI222M2R( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI222M2R$func AOI222M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI222M2R$func AOI222M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI222M4R( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI222M4R$func AOI222M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI222M4R$func AOI222M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI222M6RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI222M6RA$func AOI222M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI222M6RA$func AOI222M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI222M8RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI222M8RA$func AOI222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI222M8RA$func AOI222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22B20M0R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22B20M0R$func AOI22B20M0R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M0R$func AOI22B20M0R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22B20M1R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22B20M1R$func AOI22B20M1R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M1R$func AOI22B20M1R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22B20M2R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22B20M2R$func AOI22B20M2R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M2R$func AOI22B20M2R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22B20M4R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22B20M4R$func AOI22B20M4R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M4R$func AOI22B20M4R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22B20M8RA( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22B20M8RA$func AOI22B20M8RA_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22B20M8RA$func AOI22B20M8RA_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M0R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M0R$func AOI22M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M0R$func AOI22M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M12RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M12RA$func AOI22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M12RA$func AOI22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M16RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M16RA$func AOI22M16RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M16RA$func AOI22M16RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M1R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M1R$func AOI22M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M1R$func AOI22M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M2R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M2R$func AOI22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M2R$func AOI22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M4R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M4R$func AOI22M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M4R$func AOI22M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M6RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M6RA$func AOI22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M6RA$func AOI22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI22M8RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI22M8RA$func AOI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI22M8RA$func AOI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M0R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M0R$func AOI31M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M0R$func AOI31M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M12RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M12RA$func AOI31M12RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M12RA$func AOI31M12RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M1R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M1R$func AOI31M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M1R$func AOI31M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M2R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M2R$func AOI31M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M2R$func AOI31M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M4R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M4R$func AOI31M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M4R$func AOI31M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M6RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M6RA$func AOI31M6RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M6RA$func AOI31M6RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI31M8RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI31M8RA$func AOI31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI31M8RA$func AOI31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M0R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M0R$func AOI32M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M0R$func AOI32M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M12RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M12RA$func AOI32M12RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M12RA$func AOI32M12RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M1R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M1R$func AOI32M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M1R$func AOI32M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M2R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M2R$func AOI32M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M2R$func AOI32M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M4R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M4R$func AOI32M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M4R$func AOI32M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M6RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M6RA$func AOI32M6RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M6RA$func AOI32M6RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI32M8RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI32M8RA$func AOI32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI32M8RA$func AOI32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI33M0R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI33M0R$func AOI33M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI33M0R$func AOI33M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI33M1R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI33M1R$func AOI33M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI33M1R$func AOI33M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI33M2R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI33M2R$func AOI33M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI33M2R$func AOI33M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI33M4R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI33M4R$func AOI33M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI33M4R$func AOI33M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AOI33M8RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	AOI33M8RA$func AOI33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	AOI33M8RA$func AOI33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEM2RA( OA1, OA2, Z, M0, M1, M2);
input M0, M1, M2;
output OA1, OA2, Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEM2RA$func BEM2RA_inst(.M0(M0),.M1(M1),.M2(M2),.OA1(OA1),.OA2(OA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEM2RA$func BEM2RA_inst(.M0(M0),.M1(M1),.M2(M2),.OA1(OA1),.OA2(OA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc M0 --> OA1
	 (M0 => OA1) = (1.0,1.0);

	// arc M1 --> OA1
	 (M1 => OA1) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	ifnone
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	// arc M0 --> OA2
	 (M0 => OA2) = (1.0,1.0);

	// arc M1 --> OA2
	 (M1 => OA2) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	ifnone
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M2===1'b0)
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b0)
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b1)
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b1)
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b0)
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b0)
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b1)
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b1)
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEM4RA( OA1, OA2, Z, M0, M1, M2);
input M0, M1, M2;
output OA1, OA2, Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEM4RA$func BEM4RA_inst(.M0(M0),.M1(M1),.M2(M2),.OA1(OA1),.OA2(OA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEM4RA$func BEM4RA_inst(.M0(M0),.M1(M1),.M2(M2),.OA1(OA1),.OA2(OA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc M0 --> OA1
	 (M0 => OA1) = (1.0,1.0);

	// arc M1 --> OA1
	 (M1 => OA1) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	ifnone
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	// arc M0 --> OA2
	 (M0 => OA2) = (1.0,1.0);

	// arc M1 --> OA2
	 (M1 => OA2) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	ifnone
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M2===1'b0)
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b0)
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b1)
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b1)
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b0)
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b0)
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b1)
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b1)
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEM8RA( OA1, OA2, Z, M0, M1, M2);
input M0, M1, M2;
output OA1, OA2, Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEM8RA$func BEM8RA_inst(.M0(M0),.M1(M1),.M2(M2),.OA1(OA1),.OA2(OA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEM8RA$func BEM8RA_inst(.M0(M0),.M1(M1),.M2(M2),.OA1(OA1),.OA2(OA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc M0 --> OA1
	 (M0 => OA1) = (1.0,1.0);

	// arc M1 --> OA1
	 (M1 => OA1) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0)
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	ifnone
	// arc M2 --> OA1
	 (M2 => OA1) = (1.0,1.0);

	// arc M0 --> OA2
	 (M0 => OA2) = (1.0,1.0);

	// arc M1 --> OA2
	 (M1 => OA2) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1)
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	ifnone
	// arc M2 --> OA2
	 (M2 => OA2) = (1.0,1.0);

	if(M2===1'b0)
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b0)
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b1)
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b1)
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (Z:M0)
	 (posedge M0 => (Z:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (Z:M0)
	 (negedge M0 => (Z:M0)) = (1.0,1.0);

	if(M2===1'b0)
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b0)
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b1)
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

	if(M2===1'b1)
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (Z:M1)
	 (posedge M1 => (Z:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (Z:M1)
	 (negedge M1 => (Z:M1)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEMXBM2R( PB, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output PB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEMXBM2R$func BEMXBM2R_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.PB(PB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEMXBM2R$func BEMXBM2R_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.PB(PB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(M1===1'b0)
	// arc posedge M0 --> (PB:M0)
	 (posedge M0 => (PB:M0)) = (1.0,1.0);

	if(M1===1'b0)
	// arc negedge M0 --> (PB:M0)
	 (negedge M0 => (PB:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc posedge M0 --> (PB:M0)
	 (posedge M0 => (PB:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc negedge M0 --> (PB:M0)
	 (negedge M0 => (PB:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (PB:M0)
	 (posedge M0 => (PB:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (PB:M0)
	 (negedge M0 => (PB:M0)) = (1.0,1.0);

	if(M0===1'b0)
	// arc posedge M1 --> (PB:M1)
	 (posedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b0)
	// arc negedge M1 --> (PB:M1)
	 (negedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc posedge M1 --> (PB:M1)
	 (posedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc negedge M1 --> (PB:M1)
	 (negedge M1 => (PB:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (PB:M1)
	 (posedge M1 => (PB:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (PB:M1)
	 (negedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	ifnone
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	ifnone
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

        ifnone
	// arc posedge Z --> (PB:Z)
	 (posedge Z => (PB:Z)) = (1.0,1.0);

        ifnone
	// arc negedge Z --> (PB:Z)
	 (negedge Z => (PB:Z)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEMXBM4R( PB, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output PB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEMXBM4R$func BEMXBM4R_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.PB(PB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEMXBM4R$func BEMXBM4R_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.PB(PB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(M1===1'b0)
	// arc posedge M0 --> (PB:M0)
	 (posedge M0 => (PB:M0)) = (1.0,1.0);

	if(M1===1'b0)
	// arc negedge M0 --> (PB:M0)
	 (negedge M0 => (PB:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc posedge M0 --> (PB:M0)
	 (posedge M0 => (PB:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc negedge M0 --> (PB:M0)
	 (negedge M0 => (PB:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (PB:M0)
	 (posedge M0 => (PB:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (PB:M0)
	 (negedge M0 => (PB:M0)) = (1.0,1.0);

	if(M0===1'b0)
	// arc posedge M1 --> (PB:M1)
	 (posedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b0)
	// arc negedge M1 --> (PB:M1)
	 (negedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc posedge M1 --> (PB:M1)
	 (posedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc negedge M1 --> (PB:M1)
	 (negedge M1 => (PB:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (PB:M1)
	 (posedge M1 => (PB:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (PB:M1)
	 (negedge M1 => (PB:M1)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	ifnone
	// arc OA1 --> PB
	 (OA1 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	ifnone
	// arc OA2 --> PB
	 (OA2 => PB) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

        ifnone
	// arc posedge Z --> (PB:Z)
	 (posedge Z => (PB:Z)) = (1.0,1.0);

        ifnone
	// arc negedge Z --> (PB:Z)
	 (negedge Z => (PB:Z)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> PB
	 (Z => PB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEMXM2RA( P, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output P;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEMXM2RA$func BEMXM2RA_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.P(P),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEMXM2RA$func BEMXM2RA_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.P(P),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(M1===1'b0)
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b0)
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

	if(M0===1'b0)
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b0)
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	ifnone
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	ifnone
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

        ifnone
	// arc posedge Z --> (P:Z)
	 (posedge Z => (P:Z)) = (1.0,1.0);

        ifnone
	// arc negedge Z --> (P:Z)
	 (negedge Z => (P:Z)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEMXM4RA( P, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output P;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEMXM4RA$func BEMXM4RA_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.P(P),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEMXM4RA$func BEMXM4RA_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.P(P),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(M1===1'b0)
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b0)
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

	if(M0===1'b0)
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b0)
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	ifnone
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	ifnone
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

        ifnone
	// arc posedge Z --> (P:Z)
	 (posedge Z => (P:Z)) = (1.0,1.0);

        ifnone
	// arc negedge Z --> (P:Z)
	 (negedge Z => (P:Z)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BEMXM8RA( P, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output P;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BEMXM8RA$func BEMXM8RA_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.P(P),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BEMXM8RA$func BEMXM8RA_inst(.M0(M0),.M1(M1),.OA1(OA1),.OA2(OA2),.P(P),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(M1===1'b0)
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b0)
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

	if(M1===1'b1)
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

        ifnone
	// arc posedge M0 --> (P:M0)
	 (posedge M0 => (P:M0)) = (1.0,1.0);

        ifnone
	// arc negedge M0 --> (P:M0)
	 (negedge M0 => (P:M0)) = (1.0,1.0);

	if(M0===1'b0)
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b0)
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b1)
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

        ifnone
	// arc posedge M1 --> (P:M1)
	 (posedge M1 => (P:M1)) = (1.0,1.0);

        ifnone
	// arc negedge M1 --> (P:M1)
	 (negedge M1 => (P:M1)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	ifnone
	// arc OA1 --> P
	 (OA1 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	ifnone
	// arc OA2 --> P
	 (OA2 => P) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

        ifnone
	// arc posedge Z --> (P:Z)
	 (posedge Z => (P:Z)) = (1.0,1.0);

        ifnone
	// arc negedge Z --> (P:Z)
	 (negedge Z => (P:Z)) = (1.0,1.0);

	if(M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

	if(M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
	// arc Z --> P
	 (Z => P) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BHDM1R( Z);
inout Z;

    // Busholder.
  wire io_wire;

  buf(weak0,weak1) SMC_I0(Z, io_wire);
  buf              SMC_I1(io_wire, Z);
 
endmodule
`endcelldefine
`celldefine
module BUFM10R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM10R$func BUFM10R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM10R$func BUFM10R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM12R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM12R$func BUFM12R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM12R$func BUFM12R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM14R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM14R$func BUFM14R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM14R$func BUFM14R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM16R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM16R$func BUFM16R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM16R$func BUFM16R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM18R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM18R$func BUFM18R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM18R$func BUFM18R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM20R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM20R$func BUFM20R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM20R$func BUFM20R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM22RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM22RA$func BUFM22RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM22RA$func BUFM22RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM24R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM24R$func BUFM24R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM24R$func BUFM24R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM26RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM26RA$func BUFM26RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM26RA$func BUFM26RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM2R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM2R$func BUFM2R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM2R$func BUFM2R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM32RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM32RA$func BUFM32RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM32RA$func BUFM32RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM3R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM3R$func BUFM3R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM3R$func BUFM3R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM40RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM40RA$func BUFM40RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM40RA$func BUFM40RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM48RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM48RA$func BUFM48RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM48RA$func BUFM48RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM4R$func BUFM4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM4R$func BUFM4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM5R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM5R$func BUFM5R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM5R$func BUFM5R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM6R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM6R$func BUFM6R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM6R$func BUFM6R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFM8R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFM8R$func BUFM8R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFM8R$func BUFM8R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM0R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM0R$func BUFTM0R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM0R$func BUFTM0R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM12R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM12R$func BUFTM12R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM12R$func BUFTM12R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM16R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM16R$func BUFTM16R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM16R$func BUFTM16R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM1R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM1R$func BUFTM1R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM1R$func BUFTM1R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM20R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM20R$func BUFTM20R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM20R$func BUFTM20R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM22RA( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM22RA$func BUFTM22RA_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM22RA$func BUFTM22RA_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM24RA( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM24RA$func BUFTM24RA_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM24RA$func BUFTM24RA_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM2R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM2R$func BUFTM2R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM2R$func BUFTM2R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM32RA( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM32RA$func BUFTM32RA_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM32RA$func BUFTM32RA_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM3R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM3R$func BUFTM3R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM3R$func BUFTM3R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM40RA( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM40RA$func BUFTM40RA_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM40RA$func BUFTM40RA_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM48RA( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM48RA$func BUFTM48RA_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM48RA$func BUFTM48RA_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM4R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM4R$func BUFTM4R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM4R$func BUFTM4R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM6R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM6R$func BUFTM6R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM6R$func BUFTM6R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module BUFTM8R( Z, A, E);
input A, E;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	BUFTM8R$func BUFTM8R_inst(.A(A),.E(E),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	BUFTM8R$func BUFTM8R_inst(.A(A),.E(E),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M12R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M12R$func CKAN2M12R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M12R$func CKAN2M12R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M16RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M16RA$func CKAN2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M16RA$func CKAN2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M2R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M2R$func CKAN2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M2R$func CKAN2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M3R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M3R$func CKAN2M3R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M3R$func CKAN2M3R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M4R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M4R$func CKAN2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M4R$func CKAN2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M6R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M6R$func CKAN2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M6R$func CKAN2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKAN2M8RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKAN2M8RA$func CKAN2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKAN2M8RA$func CKAN2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM12R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM12R$func CKBUFM12R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM12R$func CKBUFM12R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM16R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM16R$func CKBUFM16R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM16R$func CKBUFM16R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM1R$func CKBUFM1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM1R$func CKBUFM1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM20R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM20R$func CKBUFM20R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM20R$func CKBUFM20R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM22RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM22RA$func CKBUFM22RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM22RA$func CKBUFM22RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM24R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM24R$func CKBUFM24R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM24R$func CKBUFM24R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM26RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM26RA$func CKBUFM26RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM26RA$func CKBUFM26RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM2R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM2R$func CKBUFM2R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM2R$func CKBUFM2R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM32R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM32R$func CKBUFM32R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM32R$func CKBUFM32R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM3R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM3R$func CKBUFM3R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM3R$func CKBUFM3R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM40R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM40R$func CKBUFM40R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM40R$func CKBUFM40R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM48R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM48R$func CKBUFM48R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM48R$func CKBUFM48R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM4R$func CKBUFM4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM4R$func CKBUFM4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM6R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM6R$func CKBUFM6R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM6R$func CKBUFM6R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKBUFM8R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKBUFM8R$func CKBUFM8R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKBUFM8R$func CKBUFM8R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM12R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM12R$func CKINVM12R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM12R$func CKINVM12R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM16R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM16R$func CKINVM16R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM16R$func CKINVM16R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM1R$func CKINVM1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM1R$func CKINVM1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM20R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM20R$func CKINVM20R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM20R$func CKINVM20R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM22RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM22RA$func CKINVM22RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM22RA$func CKINVM22RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM24R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM24R$func CKINVM24R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM24R$func CKINVM24R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM26RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM26RA$func CKINVM26RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM26RA$func CKINVM26RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM2R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM2R$func CKINVM2R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM2R$func CKINVM2R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM32R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM32R$func CKINVM32R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM32R$func CKINVM32R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM3R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM3R$func CKINVM3R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM3R$func CKINVM3R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM40R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM40R$func CKINVM40R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM40R$func CKINVM40R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM48R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM48R$func CKINVM48R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM48R$func CKINVM48R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM4R$func CKINVM4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM4R$func CKINVM4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM6R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM6R$func CKINVM6R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM6R$func CKINVM6R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKINVM8R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKINVM8R$func CKINVM8R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKINVM8R$func CKINVM8R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M12R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M12R$func CKMUX2M12R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M12R$func CKMUX2M12R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M16RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M16RA$func CKMUX2M16RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M16RA$func CKMUX2M16RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M2R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M2R$func CKMUX2M2R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M2R$func CKMUX2M2R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M3R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M3R$func CKMUX2M3R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M3R$func CKMUX2M3R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M4R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M4R$func CKMUX2M4R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M4R$func CKMUX2M4R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M6R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M6R$func CKMUX2M6R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M6R$func CKMUX2M6R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKMUX2M8R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKMUX2M8R$func CKMUX2M8R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKMUX2M8R$func CKMUX2M8R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKND2M12R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKND2M12R$func CKND2M12R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKND2M12R$func CKND2M12R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKND2M16RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKND2M16RA$func CKND2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKND2M16RA$func CKND2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKND2M2R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKND2M2R$func CKND2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKND2M2R$func CKND2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKND2M4R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKND2M4R$func CKND2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKND2M4R$func CKND2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKND2M6RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKND2M6RA$func CKND2M6RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKND2M6RA$func CKND2M6RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKND2M8R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKND2M8R$func CKND2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKND2M8R$func CKND2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKXOR2M12RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKXOR2M12RA$func CKXOR2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M12RA$func CKXOR2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKXOR2M1RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKXOR2M1RA$func CKXOR2M1RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M1RA$func CKXOR2M1RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKXOR2M2RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKXOR2M2RA$func CKXOR2M2RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M2RA$func CKXOR2M2RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKXOR2M4RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKXOR2M4RA$func CKXOR2M4RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M4RA$func CKXOR2M4RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module CKXOR2M8RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	CKXOR2M8RA$func CKXOR2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	CKXOR2M8RA$func CKXOR2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL1M1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL1M1R$func DEL1M1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL1M1R$func DEL1M1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL1M4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL1M4R$func DEL1M4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL1M4R$func DEL1M4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL2M1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL2M1R$func DEL2M1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL2M1R$func DEL2M1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL2M4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL2M4R$func DEL2M4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL2M4R$func DEL2M4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL3M1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL3M1R$func DEL3M1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL3M1R$func DEL3M1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL3M4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL3M4R$func DEL3M4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL3M4R$func DEL3M4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL4M1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL4M1R$func DEL4M1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL4M1R$func DEL4M1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DEL4M4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	DEL4M4R$func DEL4M4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DEL4M4R$func DEL4M4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFAQM1RA( Q, A, B, CK);
input A, B, CK;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;

	DFAQM1RA$func DFAQM1RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFAQM1RA$func DFAQM1RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK,negedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK,posedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,negedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,posedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFAQM2RA( Q, A, B, CK);
input A, B, CK;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;

	DFAQM2RA$func DFAQM2RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFAQM2RA$func DFAQM2RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK,negedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK,posedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,negedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,posedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFAQM4RA( Q, A, B, CK);
input A, B, CK;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;

	DFAQM4RA$func DFAQM4RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFAQM4RA$func DFAQM4RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK,negedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK,posedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,negedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,posedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFAQM6RA( Q, A, B, CK);
input A, B, CK;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;

	DFAQM6RA$func DFAQM6RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFAQM6RA$func DFAQM6RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK,negedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK,posedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,negedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,posedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFAQM8RA( Q, A, B, CK);
input A, B, CK;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;

	DFAQM8RA$func DFAQM8RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFAQM8RA$func DFAQM8RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK,negedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK,posedge A,1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,negedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK,posedge B,1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCM1RA( Q, QB, CKB, D);
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCM1RA$func DFCM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCM1RA$func DFCM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCM2RA( Q, QB, CKB, D);
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCM2RA$func DFCM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCM2RA$func DFCM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCM4RA( Q, QB, CKB, D);
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCM4RA$func DFCM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCM4RA$func DFCM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCM8RA( Q, QB, CKB, D);
input CKB, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCM8RA$func DFCM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCM8RA$func DFCM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQM1RA( Q, CKB, D);
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCQM1RA$func DFCQM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQM1RA$func DFCQM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQM2RA( Q, CKB, D);
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCQM2RA$func DFCQM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQM2RA$func DFCQM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQM4RA( Q, CKB, D);
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCQM4RA$func DFCQM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQM4RA$func DFCQM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQM8RA( Q, CKB, D);
input CKB, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;

	DFCQM8RA$func DFCQM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQM8RA$func DFCQM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,negedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB,posedge D,1.0,1.0,notifier,,,CKB$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRM1RA( Q, CKB, D, RB);
input CKB, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCQRM1RA$func DFCQRM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRM1RA$func DFCQRM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRM2RA( Q, CKB, D, RB);
input CKB, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCQRM2RA$func DFCQRM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRM2RA$func DFCQRM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRM4RA( Q, CKB, D, RB);
input CKB, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCQRM4RA$func DFCQRM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRM4RA$func DFCQRM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRM8RA( Q, CKB, D, RB);
input CKB, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCQRM8RA$func DFCQRM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRM8RA$func DFCQRM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRSM1RA( Q, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCQRSM1RA$func DFCQRSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM1RA$func DFCQRSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRSM2RA( Q, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCQRSM2RA$func DFCQRSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM2RA$func DFCQRSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRSM4RA( Q, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCQRSM4RA$func DFCQRSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM4RA$func DFCQRSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQRSM8RA( Q, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCQRSM8RA$func DFCQRSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQRSM8RA$func DFCQRSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQSM1RA( Q, CKB, D, SB);
input CKB, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCQSM1RA$func DFCQSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQSM1RA$func DFCQSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQSM2RA( Q, CKB, D, SB);
input CKB, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCQSM2RA$func DFCQSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQSM2RA$func DFCQSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQSM4RA( Q, CKB, D, SB);
input CKB, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCQSM4RA$func DFCQSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQSM4RA$func DFCQSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCQSM8RA( Q, CKB, D, SB);
input CKB, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCQSM8RA$func DFCQSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCQSM8RA$func DFCQSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRM1RA( Q, QB, CKB, D, RB);
input CKB, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCRM1RA$func DFCRM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRM1RA$func DFCRM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRM2RA( Q, QB, CKB, D, RB);
input CKB, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCRM2RA$func DFCRM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRM2RA$func DFCRM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRM4RA( Q, QB, CKB, D, RB);
input CKB, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCRM4RA$func DFCRM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRM4RA$func DFCRM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRM8RA( Q, QB, CKB, D, RB);
input CKB, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFCRM8RA$func DFCRM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRM8RA$func DFCRM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRSM1RA( Q, QB, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCRSM1RA$func DFCRSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRSM1RA$func DFCRSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRSM2RA( Q, QB, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCRSM2RA$func DFCRSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRSM2RA$func DFCRSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRSM4RA( Q, QB, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCRSM4RA$func DFCRSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRSM4RA$func DFCRSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCRSM8RA( Q, QB, CKB, D, RB, SB);
input CKB, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFCRSM8RA$func DFCRSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCRSM8RA$func DFCRSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCSM1RA( Q, QB, CKB, D, SB);
input CKB, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCSM1RA$func DFCSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCSM1RA$func DFCSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCSM2RA( Q, QB, CKB, D, SB);
input CKB, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCSM2RA$func DFCSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCSM2RA$func DFCSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCSM4RA( Q, QB, CKB, D, SB);
input CKB, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCSM4RA$func DFCSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCSM4RA$func DFCSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFCSM8RA( Q, QB, CKB, D, SB);
input CKB, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFCSM8RA$func DFCSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFCSM8RA$func DFCSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEM1RA( Q, QB, CK, D, E);
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEM1RA$func DFEM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEM1RA$func DFEM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEM2RA( Q, QB, CK, D, E);
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEM2RA$func DFEM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEM2RA$func DFEM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEM4RA( Q, QB, CK, D, E);
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEM4RA$func DFEM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEM4RA$func DFEM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEM8RA( Q, QB, CK, D, E);
input CK, D, E;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEM8RA$func DFEM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEM8RA$func DFEM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQBM1RA( QB, CK, D, E);
input CK, D, E;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQBM1RA$func DFEQBM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQBM1RA$func DFEQBM1RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQBM2RA( QB, CK, D, E);
input CK, D, E;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQBM2RA$func DFEQBM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQBM2RA$func DFEQBM2RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQBM4RA( QB, CK, D, E);
input CK, D, E;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQBM4RA$func DFEQBM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQBM4RA$func DFEQBM4RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQBM8RA( QB, CK, D, E);
input CK, D, E;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQBM8RA$func DFEQBM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQBM8RA$func DFEQBM8RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQM0RA( Q, CK, D, E);
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQM0RA$func DFEQM0RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQM0RA$func DFEQM0RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQM1RA( Q, CK, D, E);
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQM1RA$func DFEQM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQM1RA$func DFEQM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQM2RA( Q, CK, D, E);
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQM2RA$func DFEQM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQM2RA$func DFEQM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQM4RA( Q, CK, D, E);
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQM4RA$func DFEQM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQM4RA$func DFEQM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQM8RA( Q, CK, D, E);
input CK, D, E;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;

	DFEQM8RA$func DFEQM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.notifier(notifier));


	buf MGM_G0(ENABLE_E ,E$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQM8RA$func DFEQM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		negedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E === 1'b1),
		posedge D &&& (ENABLE_E === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQRM1RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQRM1RA$func DFEQRM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQRM1RA$func DFEQRM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQRM2RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQRM2RA$func DFEQRM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQRM2RA$func DFEQRM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQRM4RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQRM4RA$func DFEQRM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQRM4RA$func DFEQRM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQRM8RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQRM8RA$func DFEQRM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQRM8RA$func DFEQRM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQZRM1RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQZRM1RA$func DFEQZRM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM1RA$func DFEQZRM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQZRM2RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQZRM2RA$func DFEQZRM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM2RA$func DFEQZRM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQZRM4RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQZRM4RA$func DFEQZRM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM4RA$func DFEQZRM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEQZRM8RA( Q, CK, D, E, RB);
input CK, D, E, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEQZRM8RA$func DFEQZRM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEQZRM8RA$func DFEQZRM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFERM1RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFERM1RA$func DFERM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);



   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFERM1RA$func DFERM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFERM2RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFERM2RA$func DFERM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);



   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFERM2RA$func DFERM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFERM4RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFERM4RA$func DFERM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);



   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFERM4RA$func DFERM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFERM8RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFERM8RA$func DFERM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);



   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFERM8RA$func DFERM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEZRM1RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEZRM1RA$func DFEZRM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEZRM1RA$func DFEZRM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEZRM2RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEZRM2RA$func DFEZRM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEZRM2RA$func DFEZRM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEZRM4RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEZRM4RA$func DFEZRM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEZRM4RA$func DFEZRM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFEZRM8RA( Q, QB, CK, D, E, RB);
input CK, D, E, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;

	DFEZRM8RA$func DFEZRM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_E_AND_RB ,RB$delay,E$delay);


	buf MGM_G1(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFEZRM8RA$func DFEZRM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge E &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFM1RA( Q, QB, CK, D);
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFM1RA$func DFM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFM1RA$func DFM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFM2RA( Q, QB, CK, D);
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFM2RA$func DFM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFM2RA$func DFM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFM4RA( Q, QB, CK, D);
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFM4RA$func DFM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFM4RA$func DFM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFM8RA( Q, QB, CK, D);
input CK, D;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFM8RA$func DFM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFM8RA$func DFM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMM1RA( Q, QB, CK, D1, D2, S);
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMM1RA$func DFMM1RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMM1RA$func DFMM1RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMM2RA( Q, QB, CK, D1, D2, S);
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMM2RA$func DFMM2RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMM2RA$func DFMM2RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMM4RA( Q, QB, CK, D1, D2, S);
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMM4RA$func DFMM4RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMM4RA$func DFMM4RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMM8RA( Q, QB, CK, D1, D2, S);
input CK, D1, D2, S;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMM8RA$func DFMM8RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMM8RA$func DFMM8RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMQM1RA( Q, CK, D1, D2, S);
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMQM1RA$func DFMQM1RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMQM1RA$func DFMQM1RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMQM2RA( Q, CK, D1, D2, S);
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMQM2RA$func DFMQM2RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMQM2RA$func DFMQM2RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMQM4RA( Q, CK, D1, D2, S);
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMQM4RA$func DFMQM4RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMQM4RA$func DFMQM4RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFMQM8RA( Q, CK, D1, D2, S);
input CK, D1, D2, S;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;

	DFMQM8RA$func DFMQM8RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_S ,S$delay);


	not MGM_G1(ENABLE_NOT_S ,S$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFMQM8RA$func DFMQM8RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		negedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S === 1'b1),
		posedge D1 &&& (ENABLE_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,negedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK,posedge S,1.0,1.0,notifier,,,CK$delay,S$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBM1RA( QB, CK, D);
input CK, D;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQBM1RA$func DFQBM1RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBM1RA$func DFQBM1RA_inst(.CK(CK),.D(D),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBM2RA( QB, CK, D);
input CK, D;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQBM2RA$func DFQBM2RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBM2RA$func DFQBM2RA_inst(.CK(CK),.D(D),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBM4RA( QB, CK, D);
input CK, D;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQBM4RA$func DFQBM4RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBM4RA$func DFQBM4RA_inst(.CK(CK),.D(D),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBM8RA( QB, CK, D);
input CK, D;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQBM8RA$func DFQBM8RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBM8RA$func DFQBM8RA_inst(.CK(CK),.D(D),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBRM1RA( QB, CK, D, RB);
input CK, D, RB;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQBRM1RA$func DFQBRM1RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBRM1RA$func DFQBRM1RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBRM2RA( QB, CK, D, RB);
input CK, D, RB;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQBRM2RA$func DFQBRM2RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBRM2RA$func DFQBRM2RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBRM4RA( QB, CK, D, RB);
input CK, D, RB;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQBRM4RA$func DFQBRM4RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBRM4RA$func DFQBRM4RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQBRM8RA( QB, CK, D, RB);
input CK, D, RB;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQBRM8RA$func DFQBRM8RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQBRM8RA$func DFQBRM8RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQM1RA( Q, CK, D);
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQM1RA$func DFQM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQM1RA$func DFQM1RA_inst(.CK(CK),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQM2RA( Q, CK, D);
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQM2RA$func DFQM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQM2RA$func DFQM2RA_inst(.CK(CK),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQM4RA( Q, CK, D);
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQM4RA$func DFQM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQM4RA$func DFQM4RA_inst(.CK(CK),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQM8RA( Q, CK, D);
input CK, D;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;

	DFQM8RA$func DFQM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQM8RA$func DFQM8RA_inst(.CK(CK),.D(D),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK,negedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK,posedge D,1.0,1.0,notifier,,,CK$delay,D$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRM1RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQRM1RA$func DFQRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRM1RA$func DFQRM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRM2RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQRM2RA$func DFQRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRM2RA$func DFQRM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRM4RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQRM4RA$func DFQRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRM4RA$func DFQRM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRM8RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQRM8RA$func DFQRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRM8RA$func DFQRM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRSM1RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQRSM1RA$func DFQRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRSM1RA$func DFQRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRSM2RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQRSM2RA$func DFQRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRSM2RA$func DFQRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRSM4RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQRSM4RA$func DFQRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRSM4RA$func DFQRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQRSM8RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQRSM8RA$func DFQRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQRSM8RA$func DFQRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQSM1RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQSM1RA$func DFQSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQSM1RA$func DFQSM1RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQSM2RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQSM2RA$func DFQSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQSM2RA$func DFQSM2RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQSM4RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQSM4RA$func DFQSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQSM4RA$func DFQSM4RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQSM8RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQSM8RA$func DFQSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQSM8RA$func DFQSM8RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRM1RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQZRM1RA$func DFQZRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRM1RA$func DFQZRM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRM2RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQZRM2RA$func DFQZRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRM2RA$func DFQZRM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRM4RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQZRM4RA$func DFQZRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRM4RA$func DFQZRM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRM8RA( Q, CK, D, RB);
input CK, D, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFQZRM8RA$func DFQZRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRM8RA$func DFQZRM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRSM1RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQZRSM1RA$func DFQZRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);



  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRSM1RA$func DFQZRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRSM2RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQZRSM2RA$func DFQZRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);



  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRSM2RA$func DFQZRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRSM4RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQZRSM4RA$func DFQZRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);



  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRSM4RA$func DFQZRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZRSM8RA( Q, CK, D, RB, SB);
input CK, D, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFQZRSM8RA$func DFQZRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);



  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZRSM8RA$func DFQZRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZSM1RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQZSM1RA$func DFQZSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));
  	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZSM1RA$func DFQZSM1RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZSM2RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQZSM2RA$func DFQZSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));
  	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZSM2RA$func DFQZSM2RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZSM4RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQZSM4RA$func DFQZSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));
  	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZSM4RA$func DFQZSM4RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFQZSM8RA( Q, CK, D, SB);
input CK, D, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFQZSM8RA$func DFQZSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));
  	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFQZSM8RA$func DFQZSM8RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRM1RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFRM1RA$func DFRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRM1RA$func DFRM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRM2RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFRM2RA$func DFRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRM2RA$func DFRM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRM4RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFRM4RA$func DFRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRM4RA$func DFRM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRM8RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFRM8RA$func DFRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRM8RA$func DFRM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRSM1RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFRSM1RA$func DFRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRSM1RA$func DFRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRSM2RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFRSM2RA$func DFRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRSM2RA$func DFRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRSM4RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFRSM4RA$func DFRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRSM4RA$func DFRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFRSM8RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFRSM8RA$func DFRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFRSM8RA$func DFRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFSM1RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFSM1RA$func DFSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFSM1RA$func DFSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFSM2RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFSM2RA$func DFSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFSM2RA$func DFSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFSM4RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFSM4RA$func DFSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFSM4RA$func DFSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFSM8RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFSM8RA$func DFSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFSM8RA$func DFSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRM1RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFZRM1RA$func DFZRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRM1RA$func DFZRM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRM2RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFZRM2RA$func DFZRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRM2RA$func DFZRM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRM4RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFZRM4RA$func DFZRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRM4RA$func DFZRM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRM8RA( Q, QB, CK, D, RB);
input CK, D, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;

	DFZRM8RA$func DFZRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRM8RA$func DFZRM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        negedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
        posedge D &&& (ENABLE_RB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRSM1RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFZRSM1RA$func DFZRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRSM1RA$func DFZRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRSM2RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFZRSM2RA$func DFZRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRSM2RA$func DFZRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRSM4RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFZRSM4RA$func DFZRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRSM4RA$func DFZRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZRSM8RA( Q, QB, CK, D, RB, SB);
input CK, D, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;

	DFZRSM8RA$func DFZRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


  	buf MGM_G2(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZRSM8RA$func DFZRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,negedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK,posedge RB,1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZSM1RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFZSM1RA$func DFZSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZSM1RA$func DFZSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZSM2RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFZSM2RA$func DFZSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZSM2RA$func DFZSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZSM4RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFZSM4RA$func DFZSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZSM4RA$func DFZSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module DFZSM8RA( Q, QB, CK, D, SB);
input CK, D, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;

	DFZSM8RA$func DFZSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));
  buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	DFZSM8RA$func DFZSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        negedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
        posedge D &&& (ENABLE_SB === 1'b1),1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,negedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK,posedge SB,1.0,1.0,notifier,,,CK$delay,SB$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM0R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM0R$func INVM0R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM0R$func INVM0R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM10R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM10R$func INVM10R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM10R$func INVM10R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM12R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM12R$func INVM12R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM12R$func INVM12R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM14R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM14R$func INVM14R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM14R$func INVM14R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM16R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM16R$func INVM16R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM16R$func INVM16R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM18R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM18R$func INVM18R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM18R$func INVM18R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM1R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM1R$func INVM1R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM1R$func INVM1R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM20R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM20R$func INVM20R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM20R$func INVM20R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM22RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM22RA$func INVM22RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM22RA$func INVM22RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM24R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM24R$func INVM24R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM24R$func INVM24R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM26RA( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM26RA$func INVM26RA_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM26RA$func INVM26RA_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM2R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM2R$func INVM2R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM2R$func INVM2R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM32R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM32R$func INVM32R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM32R$func INVM32R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM3R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM3R$func INVM3R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM3R$func INVM3R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM40R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM40R$func INVM40R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM40R$func INVM40R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM48R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM48R$func INVM48R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM48R$func INVM48R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM4R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM4R$func INVM4R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM4R$func INVM4R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM5R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM5R$func INVM5R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM5R$func INVM5R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM6R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM6R$func INVM6R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM6R$func INVM6R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module INVM8R( Z, A);
input A;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	INVM8R$func INVM8R_inst(.A(A),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	INVM8R$func INVM8R_inst(.A(A),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACM1RA( Q, QB, D, GB);
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACM1RA$func LACM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACM1RA$func LACM1RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACM2RA( Q, QB, D, GB);
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACM2RA$func LACM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACM2RA$func LACM2RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACM4RA( Q, QB, D, GB);
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACM4RA$func LACM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACM4RA$func LACM4RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACM8RA( Q, QB, D, GB);
input D, GB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACM8RA$func LACM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACM8RA$func LACM8RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQM1RA( Q, D, GB);
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACQM1RA$func LACQM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQM1RA$func LACQM1RA_inst(.D(D),.GB(GB),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQM2RA( Q, D, GB);
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACQM2RA$func LACQM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQM2RA$func LACQM2RA_inst(.D(D),.GB(GB),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQM4RA( Q, D, GB);
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACQM4RA$func LACQM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQM4RA$func LACQM4RA_inst(.D(D),.GB(GB),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQM8RA( Q, D, GB);
input D, GB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;

	LACQM8RA$func LACQM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQM8RA$func LACQM8RA_inst(.D(D),.GB(GB),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB,negedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB,posedge D,1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRM1RA( Q, D, GB, RB);
input D, GB, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACQRM1RA$func LACQRM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRM1RA$func LACQRM1RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRM2RA( Q, D, GB, RB);
input D, GB, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACQRM2RA$func LACQRM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRM2RA$func LACQRM2RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRM4RA( Q, D, GB, RB);
input D, GB, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACQRM4RA$func LACQRM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRM4RA$func LACQRM4RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRM8RA( Q, D, GB, RB);
input D, GB, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACQRM8RA$func LACQRM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRM8RA$func LACQRM8RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRSM1RA( Q, D, GB, RB, SB);
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACQRSM1RA$func LACQRSM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRSM1RA$func LACQRSM1RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRSM2RA( Q, D, GB, RB, SB);
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACQRSM2RA$func LACQRSM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRSM2RA$func LACQRSM2RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRSM4RA( Q, D, GB, RB, SB);
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACQRSM4RA$func LACQRSM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRSM4RA$func LACQRSM4RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQRSM8RA( Q, D, GB, RB, SB);
input D, GB, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACQRSM8RA$func LACQRSM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQRSM8RA$func LACQRSM8RA_inst(.D(D),.GB(GB),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQSM1RA( Q, D, GB, SB);
input D, GB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACQSM1RA$func LACQSM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQSM1RA$func LACQSM1RA_inst(.D(D),.GB(GB),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQSM2RA( Q, D, GB, SB);
input D, GB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACQSM2RA$func LACQSM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQSM2RA$func LACQSM2RA_inst(.D(D),.GB(GB),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQSM4RA( Q, D, GB, SB);
input D, GB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACQSM4RA$func LACQSM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQSM4RA$func LACQSM4RA_inst(.D(D),.GB(GB),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACQSM8RA( Q, D, GB, SB);
input D, GB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACQSM8RA$func LACQSM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACQSM8RA$func LACQSM8RA_inst(.D(D),.GB(GB),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRM1RA( Q, QB, D, GB, RB);
input D, GB, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACRM1RA$func LACRM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRM1RA$func LACRM1RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRM2RA( Q, QB, D, GB, RB);
input D, GB, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACRM2RA$func LACRM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRM2RA$func LACRM2RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRM4RA( Q, QB, D, GB, RB);
input D, GB, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACRM4RA$func LACRM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRM4RA$func LACRM4RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRM8RA( Q, QB, D, GB, RB);
input D, GB, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;

	LACRM8RA$func LACRM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRM8RA$func LACRM8RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB,posedge GB,1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRSM1RA( Q, QB, D, GB, RB, SB);
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACRSM1RA$func LACRSM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRSM1RA$func LACRSM1RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRSM2RA( Q, QB, D, GB, RB, SB);
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACRSM2RA$func LACRSM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRSM2RA$func LACRSM2RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRSM4RA( Q, QB, D, GB, RB, SB);
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACRSM4RA$func LACRSM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRSM4RA$func LACRSM4RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACRSM8RA( Q, QB, D, GB, RB, SB);
input D, GB, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LACRSM8RA$func LACRSM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	buf MGM_G3(ENABLE_GB ,GB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACRSM8RA$func LACRSM8RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem RB-GB-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge GB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,GB$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge GB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,GB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_GB === 1'b1),
		posedge RB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_GB === 1'b1),
		posedge SB &&& (ENABLE_GB === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACSM1RA( Q, QB, D, GB, SB);
input D, GB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACSM1RA$func LACSM1RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACSM1RA$func LACSM1RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACSM2RA( Q, QB, D, GB, SB);
input D, GB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACSM2RA$func LACSM2RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACSM2RA$func LACSM2RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACSM4RA( Q, QB, D, GB, SB);
input D, GB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACSM4RA$func LACSM4RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACSM4RA$func LACSM4RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LACSM8RA( Q, QB, D, GB, SB);
input D, GB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire GB$delay ;
	wire SB$delay ;

	LACSM8RA$func LACSM8RA_inst(.D(D$delay),.GB(GB$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LACSM8RA$func LACSM8RA_inst(.D(D),.GB(GB),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc GB --> Q
	(negedge GB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc GB --> QB
	(negedge GB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	// setuphold D- GB-LH
	$setuphold(posedge GB &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,GB$delay,D$delay);

	$width(negedge GB,1.0,0,notifier);

	// recrem SB-GB-posedge
	$recrem(posedge SB,posedge GB,1.0,1.0,notifier,,,SB$delay,GB$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM12RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM12RA$func LAGCECSM12RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM12RA$func LAGCECSM12RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM16RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM16RA$func LAGCECSM16RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM16RA$func LAGCECSM16RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM24RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM24RA$func LAGCECSM24RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM24RA$func LAGCECSM24RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	  (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM2RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM2RA$func LAGCECSM2RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM2RA$func LAGCECSM2RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM32RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM32RA$func LAGCECSM32RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM32RA$func LAGCECSM32RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM40RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM40RA$func LAGCECSM40RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM40RA$func LAGCECSM40RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM48RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM48RA$func LAGCECSM48RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM48RA$func LAGCECSM48RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM4RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM4RA$func LAGCECSM4RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM4RA$func LAGCECSM4RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM6RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM6RA$func LAGCECSM6RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM6RA$func LAGCECSM6RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCECSM8RA( GCK, CKB, E, SE);
input CKB, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCECSM8RA$func LAGCECSM8RA_inst(.CKB(CKB$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCECSM8RA$func LAGCECSM8RA_inst(.CKB(CKB),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	ifnone
	// arc CKB --> GCK
	 (CKB => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CKB --> GCK
	 (posedge CKB => (GCK : E))  = (1.0,1.0);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold E- CKB-HL
	$setuphold(negedge CKB,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CKB$delay,E$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM12R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM12R$func LAGCEM12R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM12R$func LAGCEM12R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM16R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM16R$func LAGCEM16R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM16R$func LAGCEM16R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM20R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM20R$func LAGCEM20R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM20R$func LAGCEM20R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM2R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM2R$func LAGCEM2R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM2R$func LAGCEM2R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM3R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM3R$func LAGCEM3R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM3R$func LAGCEM3R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM4R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM4R$func LAGCEM4R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM4R$func LAGCEM4R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM6R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM6R$func LAGCEM6R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM6R$func LAGCEM6R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEM8R( GCK, CK, E);
input CK, E;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEM8R$func LAGCEM8R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEM8R$func LAGCEM8R_inst(.CK(CK),.E(E),.GCK(GCK),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b1)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM12R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM12R$func LAGCEPM12R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM12R$func LAGCEPM12R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM16R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM16R$func LAGCEPM16R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM16R$func LAGCEPM16R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM20R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM20R$func LAGCEPM20R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM20R$func LAGCEPM20R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM2R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM2R$func LAGCEPM2R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM2R$func LAGCEPM2R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM3R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM3R$func LAGCEPM3R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM3R$func LAGCEPM3R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM4R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM4R$func LAGCEPM4R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM4R$func LAGCEPM4R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM6R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM6R$func LAGCEPM6R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM6R$func LAGCEPM6R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPM8R( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPM8R$func LAGCEPM8R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPM8R$func LAGCEPM8R_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM12R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM12R$func LAGCEPOM12R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM12R$func LAGCEPOM12R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM16R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM16R$func LAGCEPOM16R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM16R$func LAGCEPOM16R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM20R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM20R$func LAGCEPOM20R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM20R$func LAGCEPOM20R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM2R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM2R$func LAGCEPOM2R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM2R$func LAGCEPOM2R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM3R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM3R$func LAGCEPOM3R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM3R$func LAGCEPOM3R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM4R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM4R$func LAGCEPOM4R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM4R$func LAGCEPOM4R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM6R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM6R$func LAGCEPOM6R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM6R$func LAGCEPOM6R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCEPOM8R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;

	LAGCEPOM8R$func LAGCEPOM8R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCEPOM8R$func LAGCEPOM8R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	(negedge CK => (GCK : E))  = (1.0,1.0);

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	(CK => GCK)  = (1.0,1.0);

	if(E===1'b0)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	if(E===1'b1)
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	ifnone
	// arc SE --> GCK
	 (SE => GCK) = (1.0,1.0);

	// arc CK --> OBS
	(negedge CK => (OBS : E))  = (1.0,1.0);

	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E,1.0,1.0,notifier,,,CK$delay,E$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM12RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM12RA$func LAGCESM12RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM12RA$func LAGCESM12RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM16RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM16RA$func LAGCESM16RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM16RA$func LAGCESM16RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM24RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM24RA$func LAGCESM24RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM24RA$func LAGCESM24RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM2RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM2RA$func LAGCESM2RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM2RA$func LAGCESM2RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM32RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM32RA$func LAGCESM32RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM32RA$func LAGCESM32RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM40RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM40RA$func LAGCESM40RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM40RA$func LAGCESM40RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM48RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM48RA$func LAGCESM48RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM48RA$func LAGCESM48RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM4RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM4RA$func LAGCESM4RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM4RA$func LAGCESM4RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM6RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM6RA$func LAGCESM6RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM6RA$func LAGCESM6RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESM8RA( GCK, CK, E, SE);
input CK, E, SE;
output GCK;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESM8RA$func LAGCESM8RA_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESM8RA$func LAGCESM8RA_inst(.CK(CK),.E(E),.GCK(GCK),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM12R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM12R$func LAGCESOM12R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM12R$func LAGCESOM12R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM16R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM16R$func LAGCESOM16R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM16R$func LAGCESOM16R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM20R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM20R$func LAGCESOM20R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM20R$func LAGCESOM20R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM2R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM2R$func LAGCESOM2R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM2R$func LAGCESOM2R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM3R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM3R$func LAGCESOM3R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM3R$func LAGCESOM3R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM4R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM4R$func LAGCESOM4R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM4R$func LAGCESOM4R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM6R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM6R$func LAGCESOM6R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM6R$func LAGCESOM6R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAGCESOM8R( GCK, OBS, CK, E, SE);
input CK, E, SE;
output GCK, OBS;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire E$delay ;
	wire SE$delay ;

	LAGCESOM8R$func LAGCESOM8R_inst(.CK(CK$delay),.E(E$delay),.GCK(GCK),.OBS(OBS),.SE(SE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAGCESOM8R$func LAGCESOM8R_inst(.CK(CK),.E(E),.GCK(GCK),.OBS(OBS),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(E===1'b0 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b0)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b1 && SE===1'b1)
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	ifnone
	// arc CK --> GCK
	 (CK => GCK) = (1.0,1.0);

	if(E===1'b0 && SE===1'b0)
	// arc CK --> GCK
	 (negedge CK => (GCK : E))  = (1.0,1.0);

	if(CK===1'b0 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b0 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b0)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	if(CK===1'b1 && SE===1'b1)
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	ifnone
	// arc E --> OBS
	 (E => OBS) = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	// setuphold E- CK-LH
	$setuphold(posedge CK,negedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK,posedge E &&& (SE === 1'b0),1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE &&& (E === 1'b0),1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAM1RA( Q, QB, D, G);
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAM1RA$func LAM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAM1RA$func LAM1RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAM2RA( Q, QB, D, G);
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAM2RA$func LAM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAM2RA$func LAM2RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAM4RA( Q, QB, D, G);
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAM4RA$func LAM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAM4RA$func LAM4RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAM8RA( Q, QB, D, G);
input D, G;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAM8RA$func LAM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAM8RA$func LAM8RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQM1RA( Q, D, G);
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAQM1RA$func LAQM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQM1RA$func LAQM1RA_inst(.D(D),.G(G),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQM2RA( Q, D, G);
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAQM2RA$func LAQM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQM2RA$func LAQM2RA_inst(.D(D),.G(G),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQM4RA( Q, D, G);
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAQM4RA$func LAQM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQM4RA$func LAQM4RA_inst(.D(D),.G(G),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQM8RA( Q, D, G);
input D, G;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;

	LAQM8RA$func LAQM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQM8RA$func LAQM8RA_inst(.D(D),.G(G),.Q(Q),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G,negedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G,posedge D,1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRM1RA( Q, D, G, RB);
input D, G, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LAQRM1RA$func LAQRM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRM1RA$func LAQRM1RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRM2RA( Q, D, G, RB);
input D, G, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LAQRM2RA$func LAQRM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRM2RA$func LAQRM2RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRM4RA( Q, D, G, RB);
input D, G, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LAQRM4RA$func LAQRM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRM4RA$func LAQRM4RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRM8RA( Q, D, G, RB);
input D, G, RB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LAQRM8RA$func LAQRM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRM8RA$func LAQRM8RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRSM1RA( Q, D, G, RB, SB);
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LAQRSM1RA$func LAQRSM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRSM1RA$func LAQRSM1RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRSM2RA( Q, D, G, RB, SB);
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LAQRSM2RA$func LAQRSM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRSM2RA$func LAQRSM2RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRSM4RA( Q, D, G, RB, SB);
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LAQRSM4RA$func LAQRSM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRSM4RA$func LAQRSM4RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQRSM8RA( Q, D, G, RB, SB);
input D, G, RB, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LAQRSM8RA$func LAQRSM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQRSM8RA$func LAQRSM8RA_inst(.D(D),.G(G),.Q(Q),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQSM1RA( Q, D, G, SB);
input D, G, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LAQSM1RA$func LAQSM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQSM1RA$func LAQSM1RA_inst(.D(D),.G(G),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQSM2RA( Q, D, G, SB);
input D, G, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LAQSM2RA$func LAQSM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQSM2RA$func LAQSM2RA_inst(.D(D),.G(G),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQSM4RA( Q, D, G, SB);
input D, G, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LAQSM4RA$func LAQSM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQSM4RA$func LAQSM4RA_inst(.D(D),.G(G),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LAQSM8RA( Q, D, G, SB);
input D, G, SB;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LAQSM8RA$func LAQSM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LAQSM8RA$func LAQSM8RA_inst(.D(D),.G(G),.Q(Q),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARM1RA( Q, QB, D, G, RB);
input D, G, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LARM1RA$func LARM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARM1RA$func LARM1RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARM2RA( Q, QB, D, G, RB);
input D, G, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LARM2RA$func LARM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARM2RA$func LARM2RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARM4RA( Q, QB, D, G, RB);
input D, G, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LARM4RA$func LARM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARM4RA$func LARM4RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARM8RA( Q, QB, D, G, RB);
input D, G, RB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;

	LARM8RA$func LARM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARM8RA$func LARM8RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		negedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB === 1'b1),
		posedge D &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB,negedge G,1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARSM1RA( Q, QB, D, G, RB, SB);
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LARSM1RA$func LARSM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARSM1RA$func LARSM1RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARSM2RA( Q, QB, D, G, RB, SB);
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LARSM2RA$func LARSM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARSM2RA$func LARSM2RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARSM4RA( Q, QB, D, G, RB, SB);
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LARSM4RA$func LARSM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARSM4RA$func LARSM4RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LARSM8RA( Q, QB, D, G, RB, SB);
input D, G, RB, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire RB$delay ;
	wire SB$delay ;

	LARSM8RA$func LARSM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.notifier(notifier));


	and MGM_G0(ENABLE_RB_AND_SB ,SB$delay,RB$delay);


	buf MGM_G1(ENABLE_SB ,SB$delay);


	buf MGM_G2(ENABLE_RB ,RB$delay);


	not MGM_G3(ENABLE_NOT_G ,G$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LARSM8RA$func LARSM8RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem RB-G-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge G &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,G$delay);

	$width(negedge RB,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge G &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,G$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB &&& (ENABLE_NOT_G === 1'b1),
		posedge RB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB &&& (ENABLE_NOT_G === 1'b1),
		posedge SB &&& (ENABLE_NOT_G === 1'b1),1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LASM1RA( Q, QB, D, G, SB);
input D, G, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LASM1RA$func LASM1RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LASM1RA$func LASM1RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LASM2RA( Q, QB, D, G, SB);
input D, G, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LASM2RA$func LASM2RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LASM2RA$func LASM2RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LASM4RA( Q, QB, D, G, SB);
input D, G, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LASM4RA$func LASM4RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LASM4RA$func LASM4RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module LASM8RA( Q, QB, D, G, SB);
input D, G, SB;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire D$delay ;
	wire G$delay ;
	wire SB$delay ;

	LASM8RA$func LASM8RA_inst(.D(D$delay),.G(G$delay),.Q(Q),.QB(QB),.SB(SB$delay),.notifier(notifier));


	buf MGM_G0(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	LASM8RA$func LASM8RA_inst(.D(D),.G(G),.Q(Q),.QB(QB),.SB(SB),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc G --> Q
	(posedge G => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc D --> QB
	 (D => QB) = (1.0,1.0);

	// arc G --> QB
	(posedge G => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		negedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	// setuphold D- G-HL
	$setuphold(negedge G &&& (ENABLE_SB === 1'b1),
		posedge D &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,G$delay,D$delay);

	$width(posedge G,1.0,0,notifier);

	// recrem SB-G-negedge
	$recrem(posedge SB,negedge G,1.0,1.0,notifier,,,SB$delay,G$delay);

	$width(negedge SB,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAO222M1RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAO222M1RA$func MAO222M1RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAO222M1RA$func MAO222M1RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAO222M2RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAO222M2RA$func MAO222M2RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAO222M2RA$func MAO222M2RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAO222M4RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAO222M4RA$func MAO222M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAO222M4RA$func MAO222M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAO222M8RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAO222M8RA$func MAO222M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAO222M8RA$func MAO222M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI2223M1RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI2223M1RA$func MAOI2223M1RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M1RA$func MAOI2223M1RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI2223M2RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI2223M2RA$func MAOI2223M2RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M2RA$func MAOI2223M2RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI2223M4RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI2223M4RA$func MAOI2223M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M4RA$func MAOI2223M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI2223M8RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI2223M8RA$func MAOI2223M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI2223M8RA$func MAOI2223M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI222M1RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI222M1RA$func MAOI222M1RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI222M1RA$func MAOI222M1RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI222M2RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI222M2RA$func MAOI222M2RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI222M2RA$func MAOI222M2RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI222M4RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI222M4RA$func MAOI222M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI222M4RA$func MAOI222M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI222M8RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI222M8RA$func MAOI222M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI222M8RA$func MAOI222M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI22M1RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI22M1RA$func MAOI22M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI22M1RA$func MAOI22M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI22M2RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI22M2RA$func MAOI22M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI22M2RA$func MAOI22M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI22M4RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI22M4RA$func MAOI22M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI22M4RA$func MAOI22M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MAOI22M8RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MAOI22M8RA$func MAOI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MAOI22M8RA$func MAOI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MOAI22M1RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MOAI22M1RA$func MOAI22M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MOAI22M1RA$func MOAI22M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MOAI22M2RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MOAI22M2RA$func MOAI22M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MOAI22M2RA$func MOAI22M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MOAI22M4RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MOAI22M4RA$func MOAI22M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MOAI22M4RA$func MOAI22M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MOAI22M8RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MOAI22M8RA$func MOAI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MOAI22M8RA$func MOAI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M0RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M0RA$func MUX2M0RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M0RA$func MUX2M0RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M12RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M12RA$func MUX2M12RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M12RA$func MUX2M12RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M1RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M1RA$func MUX2M1RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M1RA$func MUX2M1RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M2RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M2RA$func MUX2M2RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M2RA$func MUX2M2RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M3RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M3RA$func MUX2M3RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M3RA$func MUX2M3RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M4RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M4RA$func MUX2M4RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M4RA$func MUX2M4RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M6R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M6R$func MUX2M6R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M6R$func MUX2M6R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

        ifnone
	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX2M8R( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX2M8R$func MUX2M8R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX2M8R$func MUX2M8R_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX3M0RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX3M0RA$func MUX3M0RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX3M0RA$func MUX3M0RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX3M1RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX3M1RA$func MUX3M1RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX3M1RA$func MUX3M1RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX3M2RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX3M2RA$func MUX3M2RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX3M2RA$func MUX3M2RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX3M4RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX3M4RA$func MUX3M4RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX3M4RA$func MUX3M4RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX3M8RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX3M8RA$func MUX3M8RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX3M8RA$func MUX3M8RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX4M0RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX4M0RA$func MUX4M0RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX4M0RA$func MUX4M0RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX4M1RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX4M1RA$func MUX4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX4M1RA$func MUX4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX4M2RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX4M2RA$func MUX4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX4M2RA$func MUX4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX4M4R( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX4M4R$func MUX4M4R_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX4M4R$func MUX4M4R_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MUX4M8RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MUX4M8RA$func MUX4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MUX4M8RA$func MUX4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M0RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M0RA$func MXB2M0RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M0RA$func MXB2M0RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M1RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M1RA$func MXB2M1RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M1RA$func MXB2M1RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M2RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M2RA$func MXB2M2RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M2RA$func MXB2M2RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M3RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M3RA$func MXB2M3RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M3RA$func MXB2M3RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M4RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M4RA$func MXB2M4RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M4RA$func MXB2M4RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M6RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M6RA$func MXB2M6RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M6RA$func MXB2M6RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB2M8RA( Z, A, B, S);
input A, B, S;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB2M8RA$func MXB2M8RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB2M8RA$func MXB2M8RA_inst(.A(A),.B(B),.S(S),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc posedge S --> (Z:S)
	 (posedge S => (Z:S)) = (1.0,1.0);

	// arc negedge S --> (Z:S)
	 (negedge S => (Z:S)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB3M0RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB3M0RA$func MXB3M0RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB3M0RA$func MXB3M0RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB3M1RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB3M1RA$func MXB3M1RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB3M1RA$func MXB3M1RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB3M2RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB3M2RA$func MXB3M2RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB3M2RA$func MXB3M2RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB3M4RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB3M4RA$func MXB3M4RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB3M4RA$func MXB3M4RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB3M8RA( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB3M8RA$func MXB3M8RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB3M8RA$func MXB3M8RA_inst(.A(A),.B(B),.C(C),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(C===1'b0)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b0)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

	if(C===1'b1)
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB4M0RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB4M0RA$func MXB4M0RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB4M0RA$func MXB4M0RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB4M1RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB4M1RA$func MXB4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB4M1RA$func MXB4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB4M2RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB4M2RA$func MXB4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB4M2RA$func MXB4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB4M4RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB4M4RA$func MXB4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB4M4RA$func MXB4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB4M6RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB4M6RA$func MXB4M6RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB4M6RA$func MXB4M6RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module MXB4M8RA( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	MXB4M8RA$func MXB4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	MXB4M8RA$func MXB4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.S0(S0),.S1(S1),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	ifnone
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	ifnone
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S0 --> (Z:S0)
	 (posedge S0 => (Z:S0)) = (1.0,1.0);

        ifnone
	// arc negedge S0 --> (Z:S0)
	 (negedge S0 => (Z:S0)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
	// arc S0 --> Z
	 (S0 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

        ifnone
	// arc posedge S1 --> (Z:S1)
	 (posedge S1 => (Z:S1)) = (1.0,1.0);

        ifnone
	// arc negedge S1 --> (Z:S1)
	 (negedge S1 => (Z:S1)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
	// arc S1 --> Z
	 (S1 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M0R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M0R$func ND2B1M0R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M0R$func ND2B1M0R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M12RA( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M12RA$func ND2B1M12RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M12RA$func ND2B1M12RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M16RA( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M16RA$func ND2B1M16RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M16RA$func ND2B1M16RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M1R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M1R$func ND2B1M1R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M1R$func ND2B1M1R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M2R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M2R$func ND2B1M2R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M2R$func ND2B1M2R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M4R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M4R$func ND2B1M4R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M4R$func ND2B1M4R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M6RA( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M6RA$func ND2B1M6RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M6RA$func ND2B1M6RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2B1M8R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2B1M8R$func ND2B1M8R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2B1M8R$func ND2B1M8R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M0R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M0R$func ND2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M0R$func ND2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M12RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M12RA$func ND2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M12RA$func ND2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M16RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M16RA$func ND2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M16RA$func ND2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M1R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M1R$func ND2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M1R$func ND2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M2R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M2R$func ND2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M2R$func ND2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M3R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M3R$func ND2M3R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M3R$func ND2M3R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M4R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M4R$func ND2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M4R$func ND2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M5R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M5R$func ND2M5R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M5R$func ND2M5R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M6R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M6R$func ND2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M6R$func ND2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND2M8R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND2M8R$func ND2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND2M8R$func ND2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M0R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M0R$func ND3B1M0R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M0R$func ND3B1M0R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M12RA( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M12RA$func ND3B1M12RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M12RA$func ND3B1M12RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M1R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M1R$func ND3B1M1R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M1R$func ND3B1M1R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M2R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M2R$func ND3B1M2R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M2R$func ND3B1M2R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M4R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M4R$func ND3B1M4R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M4R$func ND3B1M4R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M6RA( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M6RA$func ND3B1M6RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M6RA$func ND3B1M6RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3B1M8RA( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3B1M8RA$func ND3B1M8RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3B1M8RA$func ND3B1M8RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M0R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M0R$func ND3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M0R$func ND3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M12RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M12RA$func ND3M12RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M12RA$func ND3M12RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M16RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M16RA$func ND3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M16RA$func ND3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M1R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M1R$func ND3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M1R$func ND3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M2R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M2R$func ND3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M2R$func ND3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M3R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M3R$func ND3M3R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M3R$func ND3M3R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M4RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M4RA$func ND3M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M4RA$func ND3M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M6RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M6RA$func ND3M6RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M6RA$func ND3M6RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND3M8RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND3M8RA$func ND3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND3M8RA$func ND3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B1M0R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B1M0R$func ND4B1M0R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B1M0R$func ND4B1M0R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B1M1R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B1M1R$func ND4B1M1R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B1M1R$func ND4B1M1R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B1M2R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B1M2R$func ND4B1M2R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B1M2R$func ND4B1M2R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B1M4R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B1M4R$func ND4B1M4R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B1M4R$func ND4B1M4R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B1M6RA( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B1M6RA$func ND4B1M6RA_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B1M6RA$func ND4B1M6RA_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B1M8RA( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B1M8RA$func ND4B1M8RA_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B1M8RA$func ND4B1M8RA_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B2M0R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B2M0R$func ND4B2M0R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B2M0R$func ND4B2M0R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B2M1R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B2M1R$func ND4B2M1R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B2M1R$func ND4B2M1R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B2M2R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B2M2R$func ND4B2M2R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B2M2R$func ND4B2M2R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B2M4R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B2M4R$func ND4B2M4R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B2M4R$func ND4B2M4R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4B2M8RA( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4B2M8RA$func ND4B2M8RA_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4B2M8RA$func ND4B2M8RA_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M0R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M0R$func ND4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M0R$func ND4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M16RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M16RA$func ND4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M16RA$func ND4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M1R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M1R$func ND4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M1R$func ND4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M2R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M2R$func ND4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M2R$func ND4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M4R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M4R$func ND4M4R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M4R$func ND4M4R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M6R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M6R$func ND4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M6R$func ND4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module ND4M8R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	ND4M8R$func ND4M8R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	ND4M8R$func ND4M8R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M0R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M0R$func NR2B1M0R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M0R$func NR2B1M0R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M12RA( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M12RA$func NR2B1M12RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M12RA$func NR2B1M12RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M16RA( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M16RA$func NR2B1M16RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M16RA$func NR2B1M16RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M1R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M1R$func NR2B1M1R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M1R$func NR2B1M1R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M2R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M2R$func NR2B1M2R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M2R$func NR2B1M2R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M4R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M4R$func NR2B1M4R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M4R$func NR2B1M4R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M6RA( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M6RA$func NR2B1M6RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M6RA$func NR2B1M6RA_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2B1M8R( Z, B, NA);
input B, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2B1M8R$func NR2B1M8R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2B1M8R$func NR2B1M8R_inst(.B(B),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M0R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M0R$func NR2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M0R$func NR2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M12RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M12RA$func NR2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M12RA$func NR2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M16RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M16RA$func NR2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M16RA$func NR2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M1R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M1R$func NR2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M1R$func NR2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M2R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M2R$func NR2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M2R$func NR2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M3R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M3R$func NR2M3R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M3R$func NR2M3R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M4R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M4R$func NR2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M4R$func NR2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M5R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M5R$func NR2M5R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M5R$func NR2M5R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M6R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M6R$func NR2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M6R$func NR2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR2M8R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR2M8R$func NR2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR2M8R$func NR2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3B1M0R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3B1M0R$func NR3B1M0R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3B1M0R$func NR3B1M0R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3B1M1R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3B1M1R$func NR3B1M1R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3B1M1R$func NR3B1M1R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3B1M2R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3B1M2R$func NR3B1M2R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3B1M2R$func NR3B1M2R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3B1M4R( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3B1M4R$func NR3B1M4R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3B1M4R$func NR3B1M4R_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3B1M8RA( Z, B, C, NA);
input B, C, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3B1M8RA$func NR3B1M8RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3B1M8RA$func NR3B1M8RA_inst(.B(B),.C(C),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M0R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M0R$func NR3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M0R$func NR3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M16RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M16RA$func NR3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M16RA$func NR3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M1R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M1R$func NR3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M1R$func NR3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M2R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M2R$func NR3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M2R$func NR3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M4R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M4R$func NR3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M4R$func NR3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M6R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M6R$func NR3M6R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M6R$func NR3M6R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR3M8R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR3M8R$func NR3M8R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR3M8R$func NR3M8R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B1M0R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B1M0R$func NR4B1M0R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B1M0R$func NR4B1M0R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B1M1R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B1M1R$func NR4B1M1R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B1M1R$func NR4B1M1R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B1M2R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B1M2R$func NR4B1M2R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B1M2R$func NR4B1M2R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B1M4R( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B1M4R$func NR4B1M4R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B1M4R$func NR4B1M4R_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B1M8RA( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B1M8RA$func NR4B1M8RA_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B1M8RA$func NR4B1M8RA_inst(.B(B),.C(C),.D(D),.NA(NA),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B2M0R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B2M0R$func NR4B2M0R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B2M0R$func NR4B2M0R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B2M1R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B2M1R$func NR4B2M1R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B2M1R$func NR4B2M1R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B2M2R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B2M2R$func NR4B2M2R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B2M2R$func NR4B2M2R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B2M4R( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B2M4R$func NR4B2M4R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B2M4R$func NR4B2M4R_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4B2M8RA( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4B2M8RA$func NR4B2M8RA_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4B2M8RA$func NR4B2M8RA_inst(.C(C),.D(D),.NA(NA),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc NA --> Z
	 (NA => Z) = (1.0,1.0);

	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M0R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M0R$func NR4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M0R$func NR4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M16RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M16RA$func NR4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M16RA$func NR4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M1R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M1R$func NR4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M1R$func NR4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M2R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M2R$func NR4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M2R$func NR4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M4RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M4RA$func NR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M4RA$func NR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M6R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M6R$func NR4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M6R$func NR4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module NR4M8RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	NR4M8RA$func NR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	NR4M8RA$func NR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA211M12RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA211M12RA$func OA211M12RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA211M12RA$func OA211M12RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA211M1RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA211M1RA$func OA211M1RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA211M1RA$func OA211M1RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA211M2RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA211M2RA$func OA211M2RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA211M2RA$func OA211M2RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA211M4RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA211M4RA$func OA211M4RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA211M4RA$func OA211M4RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA211M6RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA211M6RA$func OA211M6RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA211M6RA$func OA211M6RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA211M8RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA211M8RA$func OA211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA211M8RA$func OA211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M0RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M0RA$func OA21M0RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M0RA$func OA21M0RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M12RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M12RA$func OA21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M12RA$func OA21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M16RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M16RA$func OA21M16RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M16RA$func OA21M16RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M1RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M1RA$func OA21M1RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M1RA$func OA21M1RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M2RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M2RA$func OA21M2RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M2RA$func OA21M2RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M4RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M4RA$func OA21M4RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M4RA$func OA21M4RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M6RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M6RA$func OA21M6RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M6RA$func OA21M6RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA21M8RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA21M8RA$func OA21M8RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA21M8RA$func OA21M8RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA221M1RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA221M1RA$func OA221M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA221M1RA$func OA221M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA221M2RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA221M2RA$func OA221M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA221M2RA$func OA221M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA221M4RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA221M4RA$func OA221M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA221M4RA$func OA221M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA221M8RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA221M8RA$func OA221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA221M8RA$func OA221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA222M1RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA222M1RA$func OA222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA222M1RA$func OA222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA222M2RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA222M2RA$func OA222M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA222M2RA$func OA222M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA222M4RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA222M4RA$func OA222M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA222M4RA$func OA222M4RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA222M8RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA222M8RA$func OA222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA222M8RA$func OA222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M0R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M0R$func OA22M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M0R$func OA22M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M12RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M12RA$func OA22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M12RA$func OA22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M16RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M16RA$func OA22M16RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M16RA$func OA22M16RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M1R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M1R$func OA22M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M1R$func OA22M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M2R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M2R$func OA22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M2R$func OA22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M4R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M4R$func OA22M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M4R$func OA22M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M6RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M6RA$func OA22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M6RA$func OA22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA22M8RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA22M8RA$func OA22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA22M8RA$func OA22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA31M1RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA31M1RA$func OA31M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA31M1RA$func OA31M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA31M2RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA31M2RA$func OA31M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA31M2RA$func OA31M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA31M4RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA31M4RA$func OA31M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA31M4RA$func OA31M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA31M8RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA31M8RA$func OA31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA31M8RA$func OA31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA32M1RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA32M1RA$func OA32M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA32M1RA$func OA32M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA32M2RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA32M2RA$func OA32M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA32M2RA$func OA32M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA32M4RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA32M4RA$func OA32M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA32M4RA$func OA32M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA32M8RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA32M8RA$func OA32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA32M8RA$func OA32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA33M1RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA33M1RA$func OA33M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA33M1RA$func OA33M1RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA33M2RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA33M2RA$func OA33M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA33M2RA$func OA33M2RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA33M4RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA33M4RA$func OA33M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA33M4RA$func OA33M4RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OA33M8RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OA33M8RA$func OA33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OA33M8RA$func OA33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211B100M0R( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211B100M0R$func OAI211B100M0R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M0R$func OAI211B100M0R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211B100M1R( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211B100M1R$func OAI211B100M1R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M1R$func OAI211B100M1R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211B100M2R( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211B100M2R$func OAI211B100M2R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M2R$func OAI211B100M2R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211B100M4R( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211B100M4R$func OAI211B100M4R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M4R$func OAI211B100M4R_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211B100M8RA( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211B100M8RA$func OAI211B100M8RA_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211B100M8RA$func OAI211B100M8RA_inst(.A1(A1),.B(B),.C(C),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211M0R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211M0R$func OAI211M0R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211M0R$func OAI211M0R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211M1R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211M1R$func OAI211M1R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211M1R$func OAI211M1R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211M2R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211M2R$func OAI211M2R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211M2R$func OAI211M2R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211M4R( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211M4R$func OAI211M4R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211M4R$func OAI211M4R_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211M6RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211M6RA$func OAI211M6RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211M6RA$func OAI211M6RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI211M8RA( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI211M8RA$func OAI211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI211M8RA$func OAI211M8RA_inst(.A1(A1),.A2(A2),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M0R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M0R$func OAI21B01M0R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M0R$func OAI21B01M0R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M12RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M12RA$func OAI21B01M12RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M12RA$func OAI21B01M12RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M16RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M16RA$func OAI21B01M16RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M16RA$func OAI21B01M16RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M1R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M1R$func OAI21B01M1R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M1R$func OAI21B01M1R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M2R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M2R$func OAI21B01M2R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M2R$func OAI21B01M2R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M4R( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M4R$func OAI21B01M4R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M4R$func OAI21B01M4R_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M6RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M6RA$func OAI21B01M6RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M6RA$func OAI21B01M6RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B01M8RA( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B01M8RA$func OAI21B01M8RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B01M8RA$func OAI21B01M8RA_inst(.A1(A1),.A2(A2),.NB(NB),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

	ifnone
	// arc NB --> Z
	 (NB => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M0R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M0R$func OAI21B10M0R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M0R$func OAI21B10M0R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M12RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M12RA$func OAI21B10M12RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M12RA$func OAI21B10M12RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M16RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M16RA$func OAI21B10M16RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M16RA$func OAI21B10M16RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M1R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M1R$func OAI21B10M1R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M1R$func OAI21B10M1R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M2R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M2R$func OAI21B10M2R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M2R$func OAI21B10M2R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M4R( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M4R$func OAI21B10M4R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M4R$func OAI21B10M4R_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M6RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M6RA$func OAI21B10M6RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M6RA$func OAI21B10M6RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B10M8RA( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B10M8RA$func OAI21B10M8RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B10M8RA$func OAI21B10M8RA_inst(.A1(A1),.B(B),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M0R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M0R$func OAI21B20M0R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M0R$func OAI21B20M0R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M12RA( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M12RA$func OAI21B20M12RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M12RA$func OAI21B20M12RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M1R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M1R$func OAI21B20M1R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M1R$func OAI21B20M1R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M2R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M2R$func OAI21B20M2R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M2R$func OAI21B20M2R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M4R( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M4R$func OAI21B20M4R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M4R$func OAI21B20M4R_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M6RA( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M6RA$func OAI21B20M6RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M6RA$func OAI21B20M6RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21B20M8RA( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21B20M8RA$func OAI21B20M8RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21B20M8RA$func OAI21B20M8RA_inst(.B(B),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M0R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M0R$func OAI21M0R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M0R$func OAI21M0R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M12RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M12RA$func OAI21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M12RA$func OAI21M12RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M16RA( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M16RA$func OAI21M16RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M16RA$func OAI21M16RA_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M1R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M1R$func OAI21M1R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M1R$func OAI21M1R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M2R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M2R$func OAI21M2R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M2R$func OAI21M2R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M3R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M3R$func OAI21M3R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M3R$func OAI21M3R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M4R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M4R$func OAI21M4R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M4R$func OAI21M4R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M6R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M6R$func OAI21M6R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M6R$func OAI21M6R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI21M8R( Z, A1, A2, B);
input A1, A2, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI21M8R$func OAI21M8R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI21M8R$func OAI21M8R_inst(.A1(A1),.A2(A2),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI221M0R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI221M0R$func OAI221M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI221M0R$func OAI221M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI221M1R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI221M1R$func OAI221M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI221M1R$func OAI221M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI221M2R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI221M2R$func OAI221M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI221M2R$func OAI221M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI221M4R( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI221M4R$func OAI221M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI221M4R$func OAI221M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI221M6RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI221M6RA$func OAI221M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI221M6RA$func OAI221M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI221M8RA( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI221M8RA$func OAI221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI221M8RA$func OAI221M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	ifnone
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI222M0RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI222M0RA$func OAI222M0RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI222M0RA$func OAI222M0RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI222M1RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI222M1RA$func OAI222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI222M1RA$func OAI222M1RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI222M2RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI222M2RA$func OAI222M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI222M2RA$func OAI222M2RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI222M4R( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI222M4R$func OAI222M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI222M4R$func OAI222M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI222M6RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI222M6RA$func OAI222M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI222M6RA$func OAI222M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI222M8RA( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI222M8RA$func OAI222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI222M8RA$func OAI222M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.C1(C1),.C2(C2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	ifnone
	// arc C1 --> Z
	 (C1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

	ifnone
	// arc C2 --> Z
	 (C2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B10M0R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B10M0R$func OAI22B10M0R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M0R$func OAI22B10M0R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B10M1R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B10M1R$func OAI22B10M1R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M1R$func OAI22B10M1R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B10M2R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B10M2R$func OAI22B10M2R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M2R$func OAI22B10M2R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B10M4R( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B10M4R$func OAI22B10M4R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M4R$func OAI22B10M4R_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B10M8RA( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B10M8RA$func OAI22B10M8RA_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B10M8RA$func OAI22B10M8RA_inst(.A1(A1),.B1(B1),.B2(B2),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B20M0R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B20M0R$func OAI22B20M0R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M0R$func OAI22B20M0R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B20M1R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B20M1R$func OAI22B20M1R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M1R$func OAI22B20M1R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B20M2R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B20M2R$func OAI22B20M2R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M2R$func OAI22B20M2R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B20M4R( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B20M4R$func OAI22B20M4R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M4R$func OAI22B20M4R_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22B20M8RA( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22B20M8RA$func OAI22B20M8RA_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22B20M8RA$func OAI22B20M8RA_inst(.B1(B1),.B2(B2),.NA1(NA1),.NA2(NA2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(NA1===1'b0 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b0 && NA2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(NA1===1'b1 && NA2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	ifnone
	// arc NA1 --> Z
	 (NA1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

	ifnone
	// arc NA2 --> Z
	 (NA2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M0R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M0R$func OAI22M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M0R$func OAI22M0R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M12RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M12RA$func OAI22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M12RA$func OAI22M12RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M16RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M16RA$func OAI22M16RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M16RA$func OAI22M16RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M1R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M1R$func OAI22M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M1R$func OAI22M1R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M2R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M2R$func OAI22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M2R$func OAI22M2R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M4R( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M4R$func OAI22M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M4R$func OAI22M4R_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M6RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M6RA$func OAI22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M6RA$func OAI22M6RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI22M8RA( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI22M8RA$func OAI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI22M8RA$func OAI22M8RA_inst(.A1(A1),.A2(A2),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI31M0R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI31M0R$func OAI31M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI31M0R$func OAI31M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI31M1R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI31M1R$func OAI31M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI31M1R$func OAI31M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI31M2R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI31M2R$func OAI31M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI31M2R$func OAI31M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI31M4R( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI31M4R$func OAI31M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI31M4R$func OAI31M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI31M8RA( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI31M8RA$func OAI31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI31M8RA$func OAI31M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	ifnone
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI32M0R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI32M0R$func OAI32M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI32M0R$func OAI32M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI32M1R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI32M1R$func OAI32M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI32M1R$func OAI32M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI32M2R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI32M2R$func OAI32M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI32M2R$func OAI32M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI32M4R( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI32M4R$func OAI32M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI32M4R$func OAI32M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI32M8RA( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI32M8RA$func OAI32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI32M8RA$func OAI32M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI33M0R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI33M0R$func OAI33M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI33M0R$func OAI33M0R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI33M1R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI33M1R$func OAI33M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI33M1R$func OAI33M1R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI33M2R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI33M2R$func OAI33M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI33M2R$func OAI33M2R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI33M4R( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI33M4R$func OAI33M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI33M4R$func OAI33M4R_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OAI33M8RA( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OAI33M8RA$func OAI33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OAI33M8RA$func OAI33M8RA_inst(.A1(A1),.A2(A2),.A3(A3),.B1(B1),.B2(B2),.B3(B3),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	ifnone
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	ifnone
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1 && B3===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	ifnone
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	ifnone
	// arc B1 --> Z
	 (B1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	ifnone
	// arc B2 --> Z
	 (B2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b0)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && A3===1'b1)
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

	ifnone
	// arc B3 --> Z
	 (B3 => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M0R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M0R$func OR2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M0R$func OR2M0R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M12RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M12RA$func OR2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M12RA$func OR2M12RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M16RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M16RA$func OR2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M16RA$func OR2M16RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M1R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M1R$func OR2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M1R$func OR2M1R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M22RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M22RA$func OR2M22RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M22RA$func OR2M22RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M2R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M2R$func OR2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M2R$func OR2M2R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M4R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M4R$func OR2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M4R$func OR2M4R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M6R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M6R$func OR2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M6R$func OR2M6R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR2M8R( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR2M8R$func OR2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR2M8R$func OR2M8R_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M0R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M0R$func OR3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M0R$func OR3M0R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M12RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M12RA$func OR3M12RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M12RA$func OR3M12RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M16RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M16RA$func OR3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M16RA$func OR3M16RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M1R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M1R$func OR3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M1R$func OR3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M2R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M2R$func OR3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M2R$func OR3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M4R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M4R$func OR3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M4R$func OR3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M6R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M6R$func OR3M6R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M6R$func OR3M6R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR3M8RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR3M8RA$func OR3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR3M8RA$func OR3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M0R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M0R$func OR4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M0R$func OR4M0R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M12RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M12RA$func OR4M12RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M12RA$func OR4M12RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M16RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M16RA$func OR4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M16RA$func OR4M16RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M1R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M1R$func OR4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M1R$func OR4M1R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M2R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M2R$func OR4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M2R$func OR4M2R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M4RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M4RA$func OR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M4RA$func OR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M6R( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M6R$func OR4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M6R$func OR4M6R_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR4M8RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR4M8RA$func OR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR4M8RA$func OR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR6M12RA( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR6M12RA$func OR6M12RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR6M12RA$func OR6M12RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

	// arc F --> Z
	 (F => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR6M1RA( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR6M1RA$func OR6M1RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR6M1RA$func OR6M1RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

	// arc F --> Z
	 (F => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR6M2RA( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR6M2RA$func OR6M2RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR6M2RA$func OR6M2RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

	// arc F --> Z
	 (F => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR6M4RA( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR6M4RA$func OR6M4RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR6M4RA$func OR6M4RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

	// arc F --> Z
	 (F => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR6M6RA( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR6M6RA$func OR6M6RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR6M6RA$func OR6M6RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

	// arc F --> Z
	 (F => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module OR6M8RA( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	OR6M8RA$func OR6M8RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	OR6M8RA$func OR6M8RA_inst(.A(A),.B(B),.C(C),.D(D),.E(E),.F(F),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	// arc E --> Z
	 (E => Z) = (1.0,1.0);

	// arc F --> Z
	 (F => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module REG1M1R( RQB, RD, RG, RGB, WE);
input RD, RG, RGB, WE;
output RQB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire RD$delay ;
	wire WE$delay ;

	REG1M1R$func REG1M1R_inst(.RD(RD$delay),.RG(RG),.RGB(RGB),.RQB(RQB),.WE(WE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,RGB);


	and MGM_G1(ENABLE_RG_AND_NOT_RGB ,MGM_W0,RG);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	REG1M1R$func REG1M1R_inst(.RD(RD),.RG(RG),.RGB(RGB),.RQB(RQB),.WE(WE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc RD --> RQB
	 (RD => RQB) = (1.0,1.0);

	// arc RG --> RQB
	 (RG => RQB) = (1.0,1.0);

	// arc RGB --> RQB
	 (RGB => RQB) = (1.0,1.0);

	// arc WE --> RQB
	(posedge WE => (RQB : RD))  = (1.0,1.0);

	// setuphold RD- WE-HL
	$setuphold(negedge WE &&& (ENABLE_RG_AND_NOT_RGB === 1'b1),
		negedge RD &&& (ENABLE_RG_AND_NOT_RGB === 1'b1),
		1.0,1.0,notifier,,,WE$delay,RD$delay);

	// setuphold RD- WE-HL
	$setuphold(negedge WE &&& (ENABLE_RG_AND_NOT_RGB === 1'b1),
		posedge RD &&& (ENABLE_RG_AND_NOT_RGB === 1'b1),
		1.0,1.0,notifier,,,WE$delay,RD$delay);

	$width(posedge WE,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module REG2M1R( RQ1B, RQ2B, RD, RG1, RG2, WE);
input RD, RG1, RG2, WE;
output RQ1B, RQ2B;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire RD$delay ;
	wire WE$delay ;

	REG2M1R$func REG2M1R_inst(.RD(RD$delay),.RG1(RG1),.RG2(RG2),.RQ1B(RQ1B),.RQ2B(RQ2B),.WE(WE$delay),.notifier(notifier));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	REG2M1R$func REG2M1R_inst(.RD(RD),.RG1(RG1),.RG2(RG2),.RQ1B(RQ1B),.RQ2B(RQ2B),.WE(WE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc RD --> RQ1B
	 (RD => RQ1B) = (1.0,1.0);

	// arc RG1 --> RQ1B
	 (RG1 => RQ1B) = (1.0,1.0);

	if(RG2===1'b0)
	// arc WE --> RQ1B
	(posedge WE => (RQ1B : RD))  = (1.0,1.0);

	if(RG2===1'b1)
	// arc WE --> RQ1B
	(posedge WE => (RQ1B : RD))  = (1.0,1.0);

	ifnone
	// arc WE --> RQ1B
	(posedge WE => (RQ1B : RD))  = (1.0,1.0);

	// arc RD --> RQ2B
	 (RD => RQ2B) = (1.0,1.0);

	// arc RG2 --> RQ2B
	 (RG2 => RQ2B) = (1.0,1.0);

	if(RG1===1'b0)
	// arc WE --> RQ2B
	(posedge WE => (RQ2B : RD))  = (1.0,1.0);

	if(RG1===1'b1)
	// arc WE --> RQ2B
	(posedge WE => (RQ2B : RD))  = (1.0,1.0);

	ifnone
	// arc WE --> RQ2B
	(posedge WE => (RQ2B : RD))  = (1.0,1.0);

	// setuphold RD- WE-HL
	$setuphold(negedge WE,negedge RD,1.0,1.0,notifier,,,WE$delay,RD$delay);

	// setuphold RD- WE-HL
	$setuphold(negedge WE,posedge RD,1.0,1.0,notifier,,,WE$delay,RD$delay);

	$width(posedge WE,1.0,0,notifier);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module REGKM1R( RQB, RD);
input RD;
output RQB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	REGKM1R$func REGKM1R_inst(.RD(RD),.RQB(RQB));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	REGKM1R$func REGKM1R_inst(.RD(RD),.RQB(RQB));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc RD --> RQB
	 (RD => RQB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module REGKM2R( RQB, RD);
input RD;
output RQB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	REGKM2R$func REGKM2R_inst(.RD(RD),.RQB(RQB));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	REGKM2R$func REGKM2R_inst(.RD(RD),.RQB(RQB));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc RD --> RQB
	 (RD => RQB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module REGKM4R( RQB, RD);
input RD;
output RQB;

   `ifdef FUNCTIONAL  //  functional //

   `else


	REGKM4R$func REGKM4R_inst(.RD(RD),.RQB(RQB));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	REGKM4R$func REGKM4R_inst(.RD(RD),.RQB(RQB));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc RD --> RQB
	 (RD => RQB) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFAQM1RA( Q, A, B, CK, SD, SE);
input A, B, CK, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFAQM1RA$func SDFAQM1RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	not MGM_G1(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G2(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFAQM1RA$func SDFAQM1RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFAQM2RA( Q, A, B, CK, SD, SE);
input A, B, CK, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFAQM2RA$func SDFAQM2RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	not MGM_G1(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G2(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFAQM2RA$func SDFAQM2RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFAQM4RA( Q, A, B, CK, SD, SE);
input A, B, CK, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFAQM4RA$func SDFAQM4RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	not MGM_G1(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G2(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFAQM4RA$func SDFAQM4RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFAQM6RA( Q, A, B, CK, SD, SE);
input A, B, CK, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFAQM6RA$func SDFAQM6RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	not MGM_G1(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G2(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFAQM6RA$func SDFAQM6RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFAQM8RA( Q, A, B, CK, SD, SE);
input A, B, CK, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire A$delay ;
	wire B$delay ;
	wire CK$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFAQM8RA$func SDFAQM8RA_inst(.A(A$delay),.B(B$delay),.CK(CK$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	not MGM_G1(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G2(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFAQM8RA$func SDFAQM8RA_inst(.A(A),.B(B),.CK(CK),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : A))  = (1.0,1.0);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold A- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge A &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,A$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	// setuphold B- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge B &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,B$delay);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCM1RA( Q, QB, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCM1RA$func SDFCM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCM1RA$func SDFCM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCM2RA( Q, QB, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCM2RA$func SDFCM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCM2RA$func SDFCM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCM4RA( Q, QB, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCM4RA$func SDFCM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCM4RA$func SDFCM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCM8RA( Q, QB, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCM8RA$func SDFCM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCM8RA$func SDFCM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQM1RA( Q, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQM1RA$func SDFCQM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQM1RA$func SDFCQM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQM2RA( Q, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQM2RA$func SDFCQM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQM2RA$func SDFCQM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQM4RA( Q, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQM4RA$func SDFCQM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQM4RA$func SDFCQM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQM8RA( Q, CKB, D, SD, SE);
input CKB, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQM8RA$func SDFCQM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQM8RA$func SDFCQM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,negedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB,posedge SE,1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRM1RA( Q, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRM1RA$func SDFCQRM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRM1RA$func SDFCQRM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRM2RA( Q, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRM2RA$func SDFCQRM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRM2RA$func SDFCQRM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRM4RA( Q, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRM4RA$func SDFCQRM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRM4RA$func SDFCQRM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRM8RA( Q, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRM8RA$func SDFCQRM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRM8RA$func SDFCQRM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRSM1RA( Q, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRSM1RA$func SDFCQRSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM1RA$func SDFCQRSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRSM2RA( Q, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRSM2RA$func SDFCQRSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM2RA$func SDFCQRSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRSM4RA( Q, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRSM4RA$func SDFCQRSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM4RA$func SDFCQRSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQRSM8RA( Q, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQRSM8RA$func SDFCQRSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQRSM8RA$func SDFCQRSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQSM1RA( Q, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQSM1RA$func SDFCQSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQSM1RA$func SDFCQSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQSM2RA( Q, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQSM2RA$func SDFCQSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQSM2RA$func SDFCQSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQSM4RA( Q, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQSM4RA$func SDFCQSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQSM4RA$func SDFCQSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCQSM8RA( Q, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCQSM8RA$func SDFCQSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCQSM8RA$func SDFCQSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRM1RA( Q, QB, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRM1RA$func SDFCRM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRM1RA$func SDFCRM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRM2RA( Q, QB, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRM2RA$func SDFCRM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRM2RA$func SDFCRM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRM4RA( Q, QB, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRM4RA$func SDFCRM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRM4RA$func SDFCRM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRM8RA( Q, QB, CKB, D, RB, SD, SE);
input CKB, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRM8RA$func SDFCRM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRM8RA$func SDFCRM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB,negedge CKB,1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRSM1RA( Q, QB, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRSM1RA$func SDFCRSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM1RA$func SDFCRSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRSM2RA( Q, QB, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRSM2RA$func SDFCRSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM2RA$func SDFCRSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRSM4RA( Q, QB, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRSM4RA$func SDFCRSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM4RA$func SDFCRSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCRSM8RA( Q, QB, CKB, D, RB, SB, SD, SE);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCRSM8RA$func SDFCRSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCRSM8RA$func SDFCRSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem RB-CKB-negedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		negedge CKB &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CKB$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CKB-negedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		negedge CKB &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CKB$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCSM1RA( Q, QB, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCSM1RA$func SDFCSM1RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCSM1RA$func SDFCSM1RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCSM2RA( Q, QB, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCSM2RA$func SDFCSM2RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCSM2RA$func SDFCSM2RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCSM4RA( Q, QB, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCSM4RA$func SDFCSM4RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCSM4RA$func SDFCSM4RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFCSM8RA( Q, QB, CKB, D, SB, SD, SE);
input CKB, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CKB$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFCSM8RA$func SDFCSM8RA_inst(.CKB(CKB$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFCSM8RA$func SDFCSM8RA_inst(.CKB(CKB),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CKB --> Q
	(negedge CKB => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CKB --> QB
	(negedge CKB => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CKB,1.0,0,notifier);

	$width(posedge CKB,1.0,0,notifier);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// setuphold D- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,D$delay);

	// recrem SB-CKB-negedge
	$recrem(posedge SB,negedge CKB,1.0,1.0,notifier,,,SB$delay,CKB$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SD- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SD$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

	// setuphold SE- CKB-HL
	$setuphold(negedge CKB &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CKB$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEM1RA( Q, QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEM1RA$func SDFEM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEM1RA$func SDFEM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEM2RA( Q, QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEM2RA$func SDFEM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEM2RA$func SDFEM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEM4RA( Q, QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEM4RA$func SDFEM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEM4RA$func SDFEM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEM8RA( Q, QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEM8RA$func SDFEM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEM8RA$func SDFEM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQBM1RA( QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQBM1RA$func SDFEQBM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQBM1RA$func SDFEQBM1RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQBM2RA( QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQBM2RA$func SDFEQBM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQBM2RA$func SDFEQBM2RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQBM4RA( QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQBM4RA$func SDFEQBM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQBM4RA$func SDFEQBM4RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQBM8RA( QB, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQBM8RA$func SDFEQBM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQBM8RA$func SDFEQBM8RA_inst(.CK(CK),.D(D),.E(E),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQM0RA( Q, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQM0RA$func SDFEQM0RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQM0RA$func SDFEQM0RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQM1RA( Q, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQM1RA$func SDFEQM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQM1RA$func SDFEQM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQM2RA( Q, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQM2RA$func SDFEQM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQM2RA$func SDFEQM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQM4RA( Q, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQM4RA$func SDFEQM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQM4RA$func SDFEQM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQM8RA( Q, CK, D, E, SD, SE);
input CK, D, E, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQM8RA$func SDFEQM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_E_AND_NOT_SE ,MGM_W0,E$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQM8RA$func SDFEQM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQRM1RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQRM1RA$func SDFEQRM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM1RA$func SDFEQRM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQRM2RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQRM2RA$func SDFEQRM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM2RA$func SDFEQRM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQRM4RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQRM4RA$func SDFEQRM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM4RA$func SDFEQRM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQRM8RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQRM8RA$func SDFEQRM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQRM8RA$func SDFEQRM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQZRM1RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQZRM1RA$func SDFEQZRM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM1RA$func SDFEQZRM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQZRM2RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQZRM2RA$func SDFEQZRM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM2RA$func SDFEQZRM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQZRM4RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQZRM4RA$func SDFEQZRM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM4RA$func SDFEQZRM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEQZRM8RA( Q, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEQZRM8RA$func SDFEQZRM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEQZRM8RA$func SDFEQZRM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFERM1RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFERM1RA$func SDFERM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);

	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFERM1RA$func SDFERM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFERM2RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFERM2RA$func SDFERM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);

	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFERM2RA$func SDFERM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFERM4RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFERM4RA$func SDFERM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);

	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFERM4RA$func SDFERM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFERM8RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFERM8RA$func SDFERM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);

	and MGM_G6(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G7(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFERM8RA$func SDFERM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEZRM1RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEZRM1RA$func SDFEZRM1RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM1RA$func SDFEZRM1RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEZRM2RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEZRM2RA$func SDFEZRM2RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM2RA$func SDFEZRM2RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEZRM4RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEZRM4RA$func SDFEZRM4RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM4RA$func SDFEZRM4RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFEZRM8RA( Q, QB, CK, D, E, RB, SD, SE);
input CK, D, E, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire E$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFEZRM8RA$func SDFEZRM8RA_inst(.CK(CK$delay),.D(D$delay),.E(E$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,RB$delay,E$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_E_AND_RB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFEZRM8RA$func SDFEZRM8RA_inst(.CK(CK),.D(D),.E(E),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_E_AND_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold E- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge E &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,E$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFM1RA( Q, QB, CK, D, SD, SE);
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFM1RA$func SDFM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFM1RA$func SDFM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFM2RA( Q, QB, CK, D, SD, SE);
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFM2RA$func SDFM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFM2RA$func SDFM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFM4RA( Q, QB, CK, D, SD, SE);
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFM4RA$func SDFM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFM4RA$func SDFM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFM8RA( Q, QB, CK, D, SD, SE);
input CK, D, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFM8RA$func SDFM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFM8RA$func SDFM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMM1RA( Q, QB, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMM1RA$func SDFMM1RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMM1RA$func SDFMM1RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMM2RA( Q, QB, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMM2RA$func SDFMM2RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMM2RA$func SDFMM2RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMM4RA( Q, QB, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMM4RA$func SDFMM4RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMM4RA$func SDFMM4RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMM8RA( Q, QB, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMM8RA$func SDFMM8RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.QB(QB),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMM8RA$func SDFMM8RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.QB(QB),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMQM1RA( Q, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMQM1RA$func SDFMQM1RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMQM1RA$func SDFMQM1RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMQM2RA( Q, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMQM2RA$func SDFMQM2RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMQM2RA$func SDFMQM2RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMQM4RA( Q, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMQM4RA$func SDFMQM4RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMQM4RA$func SDFMQM4RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFMQM8RA( Q, CK, D1, D2, S, SD, SE);
input CK, D1, D2, S, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D1$delay ;
	wire D2$delay ;
	wire S$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFMQM8RA$func SDFMQM8RA_inst(.CK(CK$delay),.D1(D1$delay),.D2(D2$delay),.Q(Q),.S(S$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_S_AND_NOT_SE ,MGM_W0,S$delay);


	not MGM_G2(MGM_W1,S$delay);


	not MGM_G3(MGM_W2,SE$delay);


	and MGM_G4(ENABLE_NOT_S_AND_NOT_SE ,MGM_W2,MGM_W1);


	not MGM_G5(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFMQM8RA$func SDFMQM8RA_inst(.CK(CK),.D1(D1),.D2(D2),.Q(Q),.S(S),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D1))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		negedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D1- CK-LH
	$setuphold(posedge CK &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		posedge D1 &&& (ENABLE_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D1$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		negedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold D2- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		posedge D2 &&& (ENABLE_NOT_S_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D2$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold S- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge S &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,S$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBM1RA( QB, CK, D, SD, SE);
input CK, D, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBM1RA$func SDFQBM1RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBM1RA$func SDFQBM1RA_inst(.CK(CK),.D(D),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBM2RA( QB, CK, D, SD, SE);
input CK, D, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBM2RA$func SDFQBM2RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBM2RA$func SDFQBM2RA_inst(.CK(CK),.D(D),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBM4RA( QB, CK, D, SD, SE);
input CK, D, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBM4RA$func SDFQBM4RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBM4RA$func SDFQBM4RA_inst(.CK(CK),.D(D),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBM8RA( QB, CK, D, SD, SE);
input CK, D, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBM8RA$func SDFQBM8RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBM8RA$func SDFQBM8RA_inst(.CK(CK),.D(D),.QB(QB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBRM1RA( QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBRM1RA$func SDFQBRM1RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBRM1RA$func SDFQBRM1RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBRM2RA( QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBRM2RA$func SDFQBRM2RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBRM2RA$func SDFQBRM2RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBRM4RA( QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBRM4RA$func SDFQBRM4RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBRM4RA$func SDFQBRM4RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQBRM8RA( QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQBRM8RA$func SDFQBRM8RA_inst(.CK(CK$delay),.D(D$delay),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQBRM8RA$func SDFQBRM8RA_inst(.CK(CK),.D(D),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQM1RA( Q, CK, D, SD, SE);
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQM1RA$func SDFQM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQM1RA$func SDFQM1RA_inst(.CK(CK),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQM2RA( Q, CK, D, SD, SE);
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQM2RA$func SDFQM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQM2RA$func SDFQM2RA_inst(.CK(CK),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQM4RA( Q, CK, D, SD, SE);
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQM4RA$func SDFQM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQM4RA$func SDFQM4RA_inst(.CK(CK),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQM8RA( Q, CK, D, SD, SE);
input CK, D, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQM8RA$func SDFQM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(ENABLE_NOT_SE ,SE$delay);


	buf MGM_G1(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQM8RA$func SDFQM8RA_inst(.CK(CK),.D(D),.Q(Q),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRM1RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRM1RA$func SDFQRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRM1RA$func SDFQRM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRM2RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRM2RA$func SDFQRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRM2RA$func SDFQRM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRM4RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRM4RA$func SDFQRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRM4RA$func SDFQRM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRM8RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRM8RA$func SDFQRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRM8RA$func SDFQRM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRSM1RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRSM1RA$func SDFQRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM1RA$func SDFQRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRSM2RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRSM2RA$func SDFQRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM2RA$func SDFQRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRSM4RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRSM4RA$func SDFQRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM4RA$func SDFQRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQRSM8RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQRSM8RA$func SDFQRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQRSM8RA$func SDFQRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQSM1RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQSM1RA$func SDFQSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQSM1RA$func SDFQSM1RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQSM2RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQSM2RA$func SDFQSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQSM2RA$func SDFQSM2RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQSM4RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQSM4RA$func SDFQSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQSM4RA$func SDFQSM4RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQSM8RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQSM8RA$func SDFQSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQSM8RA$func SDFQSM8RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRM1RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRM1RA$func SDFQZRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G4(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM1RA$func SDFQZRM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRM2RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRM2RA$func SDFQZRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G4(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM2RA$func SDFQZRM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRM4RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRM4RA$func SDFQZRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G4(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM4RA$func SDFQZRM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRM8RA( Q, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRM8RA$func SDFQZRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G4(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRM8RA$func SDFQZRM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRSM1RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRSM1RA$func SDFQZRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);

	not MGM_G3(ENABLE_NOT_SE,SE$delay);
	not MGM_G5(MGM_W3,SE$delay);

  	and MGM_G6(ENABLE_RB_AND_NOT_SE ,MGM_W3,RB$delay);

  	buf MGM_G7(ENABLE_SE ,SE$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRSM1RA$func SDFQZRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRSM2RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRSM2RA$func SDFQZRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);

	not MGM_G3(ENABLE_NOT_SE,SE$delay);
	not MGM_G5(MGM_W3,SE$delay);

  	and MGM_G6(ENABLE_RB_AND_NOT_SE ,MGM_W3,RB$delay);

  	buf MGM_G7(ENABLE_SE ,SE$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRSM2RA$func SDFQZRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRSM4RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRSM4RA$func SDFQZRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);

	not MGM_G3(ENABLE_NOT_SE,SE$delay);
	not MGM_G5(MGM_W3,SE$delay);

  	and MGM_G6(ENABLE_RB_AND_NOT_SE ,MGM_W3,RB$delay);

  	buf MGM_G7(ENABLE_SE ,SE$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRSM4RA$func SDFQZRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZRSM8RA( Q, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZRSM8RA$func SDFQZRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);

	not MGM_G3(ENABLE_NOT_SE,SE$delay);
	not MGM_G5(MGM_W3,SE$delay);

  	and MGM_G6(ENABLE_RB_AND_NOT_SE ,MGM_W3,RB$delay);

  	buf MGM_G7(ENABLE_SE ,SE$delay);


   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZRSM8RA$func SDFQZRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZSM1RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZSM1RA$func SDFQZSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G3(ENABLE_SE ,SE$delay);

  	and MGM_G5(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZSM1RA$func SDFQZSM1RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZSM2RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZSM2RA$func SDFQZSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G3(ENABLE_SE ,SE$delay);

  	and MGM_G5(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZSM2RA$func SDFQZSM2RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZSM4RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZSM4RA$func SDFQZSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G3(ENABLE_SE ,SE$delay);

  	and MGM_G5(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZSM4RA$func SDFQZSM4RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFQZSM8RA( Q, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFQZSM8RA$func SDFQZSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

  	buf MGM_G3(ENABLE_SE ,SE$delay);

  	and MGM_G5(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFQZSM8RA$func SDFQZSM8RA_inst(.CK(CK),.D(D),.Q(Q),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRM1RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRM1RA$func SDFRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRM1RA$func SDFRM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRM2RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRM2RA$func SDFRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRM2RA$func SDFRM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRM4RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRM4RA$func SDFRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRM4RA$func SDFRM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRM8RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRM8RA$func SDFRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	and MGM_G2(ENABLE_RB_AND_SE ,SE$delay,RB$delay);


	buf MGM_G3(ENABLE_RB ,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRM8RA$func SDFRM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB,posedge CK,1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		negedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB === 1'b1),
		posedge SE &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRSM1RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRSM1RA$func SDFRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRSM1RA$func SDFRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRSM2RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRSM2RA$func SDFRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRSM2RA$func SDFRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRSM4RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRSM4RA$func SDFRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRSM4RA$func SDFRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFRSM8RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFRSM8RA$func SDFRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	buf MGM_G3(ENABLE_SB ,SB$delay);


	buf MGM_G4(ENABLE_RB ,RB$delay);


	and MGM_G5(MGM_W2,SB$delay,RB$delay);


	and MGM_G6(ENABLE_RB_AND_SB_AND_SE ,SE$delay,MGM_W2);


	and MGM_G7(ENABLE_RB_AND_SB ,SB$delay,RB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFRSM8RA$func SDFRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc RB --> Q
	(RB => Q)  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc RB --> QB
	(RB => QB)  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem RB-CK-posedge
	$recrem(posedge RB &&& (ENABLE_SB === 1'b1),
		posedge CK &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,RB$delay,CK$delay);

	$width(negedge RB,1.0,0,notifier);

	// setup RB-LH SB-LH
	$setup(posedge RB,posedge SB,1.0,notifier);

	// hold RB-LH SB-LH
	$hold(posedge SB,posedge RB,1.0,notifier);

	// recrem SB-CK-posedge
	$recrem(posedge SB &&& (ENABLE_RB === 1'b1),
		posedge CK &&& (ENABLE_RB === 1'b1),
		1.0,1.0,notifier,,,SB$delay,CK$delay);

	// setup SB-LH RB-LH
	$setup(posedge SB,posedge RB,1.0,notifier);

	// hold SB-LH RB-LH
	$hold(posedge RB,posedge SB,1.0,notifier);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_RB_AND_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		negedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB === 1'b1),
		posedge SE &&& (ENABLE_RB_AND_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFSM1RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFSM1RA$func SDFSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFSM1RA$func SDFSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFSM2RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFSM2RA$func SDFSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFSM2RA$func SDFSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFSM4RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFSM4RA$func SDFSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFSM4RA$func SDFSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFSM8RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFSM8RA$func SDFSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);


	and MGM_G2(ENABLE_SB_AND_SE ,SE$delay,SB$delay);


	buf MGM_G3(ENABLE_SB ,SB$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFSM8RA$func SDFSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc SB --> Q
	(SB => Q)  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	// arc SB --> QB
	(SB => QB)  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// recrem SB-CK-posedge
	$recrem(posedge SB,posedge CK,1.0,1.0,notifier,,,SB$delay,CK$delay);

	$width(negedge SB,1.0,0,notifier);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		negedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_SE === 1'b1),
		posedge SD &&& (ENABLE_SB_AND_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		negedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB === 1'b1),
		posedge SE &&& (ENABLE_SB === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRM1RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRM1RA$func SDFZRM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRM1RA$func SDFZRM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRM2RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRM2RA$func SDFZRM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRM2RA$func SDFZRM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRM4RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRM4RA$func SDFZRM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRM4RA$func SDFZRM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRM8RA( Q, QB, CK, D, RB, SD, SE);
input CK, D, RB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRM8RA$func SDFZRM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_RB_AND_NOT_SE ,MGM_W0,RB$delay);


	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRM8RA$func SDFZRM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRSM1RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRSM1RA$func SDFZRSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(ENABLE_NOT_SE ,SE$delay);


	not MGM_G4(MGM_W2,SE$delay);


	and MGM_G5(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRSM1RA$func SDFZRSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRSM2RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRSM2RA$func SDFZRSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(ENABLE_NOT_SE ,SE$delay);


	not MGM_G4(MGM_W2,SE$delay);


	and MGM_G5(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRSM2RA$func SDFZRSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRSM4RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRSM4RA$func SDFZRSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(ENABLE_NOT_SE ,SE$delay);


	not MGM_G4(MGM_W2,SE$delay);


	and MGM_G5(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRSM4RA$func SDFZRSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZRSM8RA( Q, QB, CK, D, RB, SB, SD, SE);
input CK, D, RB, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire RB$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZRSM8RA$func SDFZRSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.RB(RB$delay),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	and MGM_G0(MGM_W0,SB$delay,RB$delay);


	not MGM_G1(MGM_W1,SE$delay);


	and MGM_G2(ENABLE_RB_AND_SB_AND_NOT_SE ,MGM_W1,MGM_W0);


	not MGM_G3(ENABLE_NOT_SE ,SE$delay);


	not MGM_G4(MGM_W2,SE$delay);


	and MGM_G5(ENABLE_RB_AND_NOT_SE ,MGM_W2,RB$delay);


	buf MGM_G6(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZRSM8RA$func SDFZRSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.RB(RB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_RB_AND_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold RB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge RB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,RB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_RB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZSM1RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZSM1RA$func SDFZSM1RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZSM1RA$func SDFZSM1RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZSM2RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZSM2RA$func SDFZSM2RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZSM2RA$func SDFZSM2RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZSM4RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZSM4RA$func SDFZSM4RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZSM4RA$func SDFZSM4RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module SDFZSM8RA( Q, QB, CK, D, SB, SD, SE);
input CK, D, SB, SD, SE;
output Q, QB;
reg notifier;

   `ifdef FUNCTIONAL  //  functional //

   `else

	wire CK$delay ;
	wire D$delay ;
	wire SB$delay ;
	wire SD$delay ;
	wire SE$delay ;

	SDFZSM8RA$func SDFZSM8RA_inst(.CK(CK$delay),.D(D$delay),.Q(Q),.QB(QB),.SB(SB$delay),.SD(SD$delay),.SE(SE$delay),.notifier(notifier));


	not MGM_G0(MGM_W0,SE$delay);


	and MGM_G1(ENABLE_SB_AND_NOT_SE ,MGM_W0,SB$delay);

	not MGM_G2(ENABLE_NOT_SE ,SE$delay);

	buf MGM_G3(ENABLE_SE ,SE$delay);

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	SDFZSM8RA$func SDFZSM8RA_inst(.CK(CK),.D(D),.Q(Q),.QB(QB),.SB(SB),.SD(SD),.SE(SE),.notifier(notifier));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	// arc CK --> QB
	(posedge CK => (QB : D))  = (1.0,1.0);

	$width(negedge CK,1.0,0,notifier);

	$width(posedge CK,1.0,0,notifier);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		negedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold D- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		posedge D &&& (ENABLE_SB_AND_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,D$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		negedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SB- CK-LH
	$setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1),
		posedge SB &&& (ENABLE_NOT_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SB$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		negedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SD- CK-LH
	$setuphold(posedge CK &&& (ENABLE_SE === 1'b1),
		posedge SD &&& (ENABLE_SE === 1'b1),
		1.0,1.0,notifier,,,CK$delay,SD$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,negedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

	// setuphold SE- CK-LH
	$setuphold(posedge CK,posedge SE,1.0,1.0,notifier,,,CK$delay,SE$delay);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module TIE0R( Z);
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	TIE0R$func TIE0R_inst(.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	TIE0R$func TIE0R_inst(.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module TIE1R( Z);
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	TIE1R$func TIE1R_inst(.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	TIE1R$func TIE1R_inst(.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR2M0RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR2M0RA$func XNR2M0RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR2M0RA$func XNR2M0RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR2M1RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR2M1RA$func XNR2M1RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR2M1RA$func XNR2M1RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR2M2RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR2M2RA$func XNR2M2RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR2M2RA$func XNR2M2RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR2M4RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR2M4RA$func XNR2M4RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR2M4RA$func XNR2M4RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR2M6RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR2M6RA$func XNR2M6RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR2M6RA$func XNR2M6RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR2M8RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR2M8RA$func XNR2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR2M8RA$func XNR2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR3M0RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR3M0RA$func XNR3M0RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR3M0RA$func XNR3M0RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR3M1R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR3M1R$func XNR3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR3M1R$func XNR3M1R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR3M2R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR3M2R$func XNR3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR3M2R$func XNR3M2R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR3M4R( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR3M4R$func XNR3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR3M4R$func XNR3M4R_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR3M6RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR3M6RA$func XNR3M6RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR3M6RA$func XNR3M6RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR3M8RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR3M8RA$func XNR3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR3M8RA$func XNR3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR4M1RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR4M1RA$func XNR4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR4M1RA$func XNR4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR4M2RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR4M2RA$func XNR4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR4M2RA$func XNR4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR4M4RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR4M4RA$func XNR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR4M4RA$func XNR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XNR4M8RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XNR4M8RA$func XNR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XNR4M8RA$func XNR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M0RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M0RA$func XOR2M0RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M0RA$func XOR2M0RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M1RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M1RA$func XOR2M1RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M1RA$func XOR2M1RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M2RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M2RA$func XOR2M2RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M2RA$func XOR2M2RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M3RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M3RA$func XOR2M3RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M3RA$func XOR2M3RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M4RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M4RA$func XOR2M4RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M4RA$func XOR2M4RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M6RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M6RA$func XOR2M6RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M6RA$func XOR2M6RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR2M8RA( Z, A, B);
input A, B;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR2M8RA$func XOR2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR2M8RA$func XOR2M8RA_inst(.A(A),.B(B),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR3M0RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR3M0RA$func XOR3M0RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR3M0RA$func XOR3M0RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR3M1RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR3M1RA$func XOR3M1RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR3M1RA$func XOR3M1RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR3M2RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR3M2RA$func XOR3M2RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR3M2RA$func XOR3M2RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR3M4RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR3M4RA$func XOR3M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR3M4RA$func XOR3M4RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR3M6RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR3M6RA$func XOR3M6RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR3M6RA$func XOR3M6RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR3M8RA( Z, A, B, C);
input A, B, C;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR3M8RA$func XOR3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR3M8RA$func XOR3M8RA_inst(.A(A),.B(B),.C(C),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR4M1RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR4M1RA$func XOR4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR4M1RA$func XOR4M1RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR4M2RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR4M2RA$func XOR4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR4M2RA$func XOR4M2RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR4M4RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR4M4RA$func XOR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR4M4RA$func XOR4M4RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module XOR4M8RA( Z, A, B, C, D);
input A, B, C, D;
output Z;

   `ifdef FUNCTIONAL  //  functional //

   `else


	XOR4M8RA$func XOR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 



   `ifdef FUNCTIONAL  //  functional //

	XOR4M8RA$func XOR4M8RA_inst(.A(A),.B(B),.C(C),.D(D),.Z(Z));

   `endif 


   `ifdef FUNCTIONAL // functional  //

   `else


// specify block begins 

   specify

	if(B===1'b0 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

        ifnone
	// arc posedge A --> (Z:A)
	 (posedge A => (Z:A)) = (1.0,1.0);

        ifnone
	// arc negedge A --> (Z:A)
	 (negedge A => (Z:A)) = (1.0,1.0);

	if(B===1'b0 && C===1'b0 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b0 && C===1'b1 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b0 && D===1'b1)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(B===1'b1 && C===1'b1 && D===1'b0)
	// arc A --> Z
	 (A => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

        ifnone
	// arc posedge B --> (Z:B)
	 (posedge B => (Z:B)) = (1.0,1.0);

        ifnone
	// arc negedge B --> (Z:B)
	 (negedge B => (Z:B)) = (1.0,1.0);

	if(A===1'b0 && C===1'b0 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && C===1'b1 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b0 && D===1'b1)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b1 && C===1'b1 && D===1'b0)
	// arc B --> Z
	 (B => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

        ifnone
	// arc posedge C --> (Z:C)
	 (posedge C => (Z:C)) = (1.0,1.0);

        ifnone
	// arc negedge C --> (Z:C)
	 (negedge C => (Z:C)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && D===1'b1)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && D===1'b0)
	// arc C --> Z
	 (C => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

        ifnone
	// arc posedge D --> (Z:D)
	 (posedge D => (Z:D)) = (1.0,1.0);

        ifnone
	// arc negedge D --> (Z:D)
	 (negedge D => (Z:D)) = (1.0,1.0);

	if(A===1'b0 && B===1'b0 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b0 && B===1'b1 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b0 && C===1'b1)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

	if(A===1'b1 && B===1'b1 && C===1'b0)
	// arc D --> Z
	 (D => Z) = (1.0,1.0);

   endspecify

   `endif 

endmodule
`endcelldefine
`celldefine
module AD42M2RA$func( CO, ICO, S, A, B, C, D, ICI);
input A, B, C, D, ICI;
output CO, ICO, S;

	AD42M2RA_udp_0(CO,A,B,C,D,ICI); 

	AD42M2RA_udp_1(ICO,A,B,C); 

	AD42M2RA_udp_2(S,A,B,C,D,ICI); 
endmodule
`endcelldefine
`celldefine
module AD42M4RA$func( CO, ICO, S, A, B, C, D, ICI);
input A, B, C, D, ICI;
output CO, ICO, S;

	AD42M2RA_udp_0(CO,A,B,C,D,ICI); 

	AD42M2RA_udp_1(ICO,A,B,C); 

	AD42M2RA_udp_2(S,A,B,C,D,ICI); 
endmodule
`endcelldefine
`celldefine
module ADCSCM2R$func( CO0, CO1, A, B, NCI0, NCI1);
input A, B, NCI0, NCI1;
output CO0, CO1;

	ADCSCM2R_udp_0(CO0,A,B,NCI0); 

	ADCSCM2R_udp_0(CO1,A,B,NCI1); 
endmodule
`endcelldefine
`celldefine
module ADCSCM4R$func( CO0, CO1, A, B, NCI0, NCI1);
input A, B, NCI0, NCI1;
output CO0, CO1;

	ADCSCM2R_udp_0(CO0,A,B,NCI0); 

	ADCSCM2R_udp_0(CO1,A,B,NCI1); 
endmodule
`endcelldefine
`celldefine
module ADCSIOM2R$func( CO0B, CO1B, A, B);
input A, B;
output CO0B, CO1B;

	ADCSIOM2R_udp_0(CO0B,A,B); 

	ADCSIOM2R_udp_1(CO1B,A,B); 
endmodule
`endcelldefine
`celldefine
module ADCSIOM4R$func( CO0B, CO1B, A, B);
input A, B;
output CO0B, CO1B;

	ADCSIOM2R_udp_0(CO0B,A,B); 

	ADCSIOM2R_udp_1(CO1B,A,B); 
endmodule
`endcelldefine
`celldefine
module ADCSOM2R$func( CO0B, CO1B, A, B, CI0, CI1);
input A, B, CI0, CI1;
output CO0B, CO1B;

	ADCSOM2R_udp_0(CO0B,A,B,CI0); 

	ADCSOM2R_udp_0(CO1B,A,B,CI1); 
endmodule
`endcelldefine
`celldefine
module ADCSOM4R$func( CO0B, CO1B, A, B, CI0, CI1);
input A, B, CI0, CI1;
output CO0B, CO1B;

	ADCSOM2R_udp_0(CO0B,A,B,CI0); 

	ADCSOM2R_udp_0(CO1B,A,B,CI1); 
endmodule
`endcelldefine
`celldefine
module ADFCGCM2RA$func( CO, A, B, NCI);
input A, B, NCI;
output CO;

	ADCSCM2R_udp_0(CO,A,B,NCI); 
endmodule
`endcelldefine
`celldefine
module ADFCGCM4RA$func( CO, A, B, NCI);
input A, B, NCI;
output CO;

	ADCSCM2R_udp_0(CO,A,B,NCI); 
endmodule
`endcelldefine
`celldefine
module ADFCGOM2RA$func( COB, A, B, CI);
input A, B, CI;
output COB;

	ADCSOM2R_udp_0(COB,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFCGOM4RA$func( COB, A, B, CI);
input A, B, CI;
output COB;

	ADCSOM2R_udp_0(COB,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFCM2RA$func( CO, S, A, B, NCI);
input A, B, NCI;
output CO, S;

	ADCSCM2R_udp_0(CO,A,B,NCI); 

	ADFCM2RA_udp_0(S,A,B,NCI); 
endmodule
`endcelldefine
`celldefine
module ADFCM4RA$func( CO, S, A, B, NCI);
input A, B, NCI;
output CO, S;

	ADCSCM2R_udp_0(CO,A,B,NCI); 

	ADFCM2RA_udp_0(S,A,B,NCI); 
endmodule
`endcelldefine
`celldefine
module ADFCSCM2RA$func( CO0, CO1, S, A, B, CS, NCI0, NCI1);
input A, B, CS, NCI0, NCI1;
output CO0, CO1, S;

	ADCSCM2R_udp_0(CO0,A,B,NCI0); 

	ADCSCM2R_udp_0(CO1,A,B,NCI1); 

	ADFCSCM2RA_udp_0(S,A,B,CS,NCI1,NCI0); 
endmodule
`endcelldefine
`celldefine
module ADFCSCM4RA$func( CO0, CO1, S, A, B, CS, NCI0, NCI1);
input A, B, CS, NCI0, NCI1;
output CO0, CO1, S;

	ADCSCM2R_udp_0(CO0,A,B,NCI0); 

	ADCSCM2R_udp_0(CO1,A,B,NCI1); 

	ADFCSCM2RA_udp_0(S,A,B,CS,NCI1,NCI0); 
endmodule
`endcelldefine
`celldefine
module ADFCSIOM2R$func( CO0B, CO1B, S, A, B, CS);
input A, B, CS;
output CO0B, CO1B, S;

	ADCSIOM2R_udp_0(CO0B,A,B); 

	ADCSIOM2R_udp_1(CO1B,A,B); 

	ADFCSIOM2R_udp_0(S,A,B,CS); 
endmodule
`endcelldefine
`celldefine
module ADFCSIOM4R$func( CO0B, CO1B, S, A, B, CS);
input A, B, CS;
output CO0B, CO1B, S;

	ADCSIOM2R_udp_0(CO0B,A,B); 

	ADCSIOM2R_udp_1(CO1B,A,B); 

	ADFCSIOM2R_udp_0(S,A,B,CS); 
endmodule
`endcelldefine
`celldefine
module ADFCSOM2RA$func( CO0B, CO1B, S, A, B, CI0, CI1, CS);
input A, B, CI0, CI1, CS;
output CO0B, CO1B, S;

	ADCSOM2R_udp_0(CO0B,A,B,CI0); 

	ADCSOM2R_udp_0(CO1B,A,B,CI1); 

	ADFCSOM2RA_udp_0(S,A,B,CI0,CS,CI1); 
endmodule
`endcelldefine
`celldefine
module ADFCSOM4RA$func( CO0B, CO1B, S, A, B, CI0, CI1, CS);
input A, B, CI0, CI1, CS;
output CO0B, CO1B, S;

	ADCSOM2R_udp_0(CO0B,A,B,CI0); 

	ADCSOM2R_udp_0(CO1B,A,B,CI1); 

	ADFCSOM2RA_udp_0(S,A,B,CI0,CS,CI1); 
endmodule
`endcelldefine
`celldefine
module ADFM0RA$func( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

	AD42M2RA_udp_1(CO,A,B,CI); 

	ADFCSIOM2R_udp_0(S,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFM1RA$func( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

	AD42M2RA_udp_1(CO,A,B,CI); 

	ADFCSIOM2R_udp_0(S,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFM2RA$func( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

	AD42M2RA_udp_1(CO,A,B,CI); 

	ADFCSIOM2R_udp_0(S,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFM4RA$func( CO, S, A, B, CI);
input A, B, CI;
output CO, S;

	AD42M2RA_udp_1(CO,A,B,CI); 

	ADFCSIOM2R_udp_0(S,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFOM2RA$func( COB, S, A, B, CI);
input A, B, CI;
output COB, S;

	ADCSOM2R_udp_0(COB,A,B,CI); 

	ADFCSIOM2R_udp_0(S,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADFOM4RA$func( COB, S, A, B, CI);
input A, B, CI;
output COB, S;

	ADCSOM2R_udp_0(COB,A,B,CI); 

	ADFCSIOM2R_udp_0(S,A,B,CI); 
endmodule
`endcelldefine
`celldefine
module ADHCM2R$func( CO, S, A, NCI);
input A, NCI;
output CO, S;

	ADHCM2R_udp_0(CO,A,NCI); 

	ADHCM2R_udp_1(S,A,NCI); 
endmodule
`endcelldefine
`celldefine
module ADHCM4R$func( CO, S, A, NCI);
input A, NCI;
output CO, S;

	ADHCM2R_udp_0(CO,A,NCI); 

	ADHCM2R_udp_1(S,A,NCI); 
endmodule
`endcelldefine
`celldefine
module ADHCSCM2R$func( CO, S, A, CS, NCI);
input A, CS, NCI;
output CO, S;

	ADHCM2R_udp_0(CO,A,NCI); 

	ADHCSCM2R_udp_0(S,A,CS,NCI); 
endmodule
`endcelldefine
`celldefine
module ADHCSCM4R$func( CO, S, A, CS, NCI);
input A, CS, NCI;
output CO, S;

	ADHCM2R_udp_0(CO,A,NCI); 

	ADHCSCM2R_udp_0(S,A,CS,NCI); 
endmodule
`endcelldefine
`celldefine
module ADHCSOM2R$func( COB, S, A, CI, CS);
input A, CI, CS;
output COB, S;

	ADCSIOM2R_udp_0(COB,A,CI); 

	ADHCSOM2R_udp_0(S,A,CI,CS); 
endmodule
`endcelldefine
`celldefine
module ADHCSOM4R$func( COB, S, A, CI, CS);
input A, CI, CS;
output COB, S;

	ADCSIOM2R_udp_0(COB,A,CI); 

	ADHCSOM2R_udp_0(S,A,CI,CS); 
endmodule
`endcelldefine
`celldefine
module ADHM1RA$func( CO, S, A, B);
input A, B;
output CO, S;

	ADHM1RA_udp_0(CO,A,B); 

	ADHM1RA_udp_1(S,A,B); 
endmodule
`endcelldefine
`celldefine
module ADHM2RA$func( CO, S, A, B);
input A, B;
output CO, S;

	ADHM1RA_udp_0(CO,A,B); 

	ADHM1RA_udp_1(S,A,B); 
endmodule
`endcelldefine
`celldefine
module ADHM4RA$func( CO, S, A, B);
input A, B;
output CO, S;

	ADHM1RA_udp_0(CO,A,B); 

	ADHM1RA_udp_1(S,A,B); 
endmodule
`endcelldefine
`celldefine
module ADHM8RA$func( CO, S, A, B);
input A, B;
output CO, S;

	ADHM1RA_udp_0(CO,A,B); 

	ADHM1RA_udp_1(S,A,B); 
endmodule
`endcelldefine
`celldefine
module ADHOM2R$func( COB, S, A, CI);
input A, CI;
output COB, S;

	ADCSIOM2R_udp_0(COB,A,CI); 

	ADHM1RA_udp_1(S,A,CI); 
endmodule
`endcelldefine
`celldefine
module ADHOM4R$func( COB, S, A, CI);
input A, CI;
output COB, S;

	ADCSIOM2R_udp_0(COB,A,CI); 

	ADHM1RA_udp_1(S,A,CI); 
endmodule
`endcelldefine
`celldefine
module AN2M0R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M12RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M16RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M1R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M22RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M2R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M4R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M6R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN2M8R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module AN3M0R$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M12RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M16RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M1R$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M22RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M2R$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M4R$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M6R$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN3M8R$func( Z, A, B, C);
input A, B, C;
output Z;

	AN3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module AN4M0R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M12RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M16RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M1R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M2R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M4RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M6R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AN4M8RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	AN4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module AO211M1RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AO211M1RA_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module AO211M2RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AO211M1RA_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module AO211M4RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AO211M1RA_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module AO211M8RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AO211M1RA_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module AO21M0RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO21M12RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO21M1RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO21M2RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO21M4RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO21M6RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO21M8RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AO21M0RA_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module AO221M1RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AO221M1RA_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module AO221M2RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AO221M1RA_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module AO221M4RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AO221M1RA_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module AO221M8RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AO221M1RA_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module AO222M1RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AO222M1RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module AO222M2RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AO222M1RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module AO222M4RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AO222M1RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module AO222M8RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AO222M1RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module AO22B10M0R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	AO22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22B10M1R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	AO22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22B10M2R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	AO22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22B10M4R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	AO22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22B10M8RA$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	AO22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22B11M0R$func( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

	AO22B11M0R_udp_0(Z,A1,NA2,B1,NB2); 
endmodule
`endcelldefine
`celldefine
module AO22B11M1R$func( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

	AO22B11M0R_udp_0(Z,A1,NA2,B1,NB2); 
endmodule
`endcelldefine
`celldefine
module AO22B11M2R$func( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

	AO22B11M0R_udp_0(Z,A1,NA2,B1,NB2); 
endmodule
`endcelldefine
`celldefine
module AO22B11M4R$func( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

	AO22B11M0R_udp_0(Z,A1,NA2,B1,NB2); 
endmodule
`endcelldefine
`celldefine
module AO22B11M8RA$func( Z, A1, B1, NA2, NB2);
input A1, B1, NA2, NB2;
output Z;

	AO22B11M0R_udp_0(Z,A1,NA2,B1,NB2); 
endmodule
`endcelldefine
`celldefine
module AO22M0RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22M12RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22M1RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22M2R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22M4RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22M6RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO22M8RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AO22M0RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO31M1RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AO31M1RA_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module AO31M2RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AO31M1RA_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module AO31M4RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AO31M1RA_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module AO31M8RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AO31M1RA_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module AO32M1RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AO32M1RA_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO32M2RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AO32M1RA_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO32M4RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AO32M1RA_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO32M8RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AO32M1RA_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module AO33M1RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AO33M1RA_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module AO33M2RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AO33M1RA_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module AO33M4RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AO33M1RA_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module AO33M8RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AO33M1RA_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module AOI211M0R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AOI211M0R_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module AOI211M1R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AOI211M0R_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module AOI211M2R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AOI211M0R_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module AOI211M4R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AOI211M0R_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module AOI211M6RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AOI211M0R_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module AOI211M8RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	AOI211M0R_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M0R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M12RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M16RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M1R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M2R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M4R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M6RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B01M8RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	AOI21B01M0R_udp_0(Z,A1,NB,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M0R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M12RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M16RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M1R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M2R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M4R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M6RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B10M8RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	AOI21B10M0R_udp_0(Z,A1,B,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B20M0R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	AOI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B20M1R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	AOI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B20M2R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	AOI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B20M4R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	AOI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21B20M8RA$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	AOI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module AOI21M0R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M12RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M16RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M1R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M2R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M3R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M4R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M6R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI21M8R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	AOI21M0R_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module AOI221M0R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AOI221M0R_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI221M1R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AOI221M0R_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI221M2R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AOI221M0R_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI221M4R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AOI221M0R_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI221M6RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AOI221M0R_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI221M8RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	AOI221M0R_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI222M0RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AOI222M0RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI222M1RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AOI222M0RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI222M2R$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AOI222M0RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI222M4R$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AOI222M0RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI222M6RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AOI222M0RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI222M8RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	AOI222M0RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22B20M0R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	AOI22B20M0R_udp_0(Z,B1,NA1,NA2,B2); 
endmodule
`endcelldefine
`celldefine
module AOI22B20M1R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	AOI22B20M0R_udp_0(Z,B1,NA1,NA2,B2); 
endmodule
`endcelldefine
`celldefine
module AOI22B20M2R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	AOI22B20M0R_udp_0(Z,B1,NA1,NA2,B2); 
endmodule
`endcelldefine
`celldefine
module AOI22B20M4R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	AOI22B20M0R_udp_0(Z,B1,NA1,NA2,B2); 
endmodule
`endcelldefine
`celldefine
module AOI22B20M8RA$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	AOI22B20M0R_udp_0(Z,B1,NA1,NA2,B2); 
endmodule
`endcelldefine
`celldefine
module AOI22M0R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M12RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M16RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M1R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M2R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M4R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M6RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI22M8RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module AOI31M0R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI31M12RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI31M1R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI31M2R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI31M4R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI31M6RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI31M8RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	AOI31M0R_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M0R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M12RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M1R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M2R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M4R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M6RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI32M8RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	AOI32M0R_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI33M0R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AOI33M0R_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI33M1R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AOI33M0R_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI33M2R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AOI33M0R_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI33M4R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AOI33M0R_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module AOI33M8RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	AOI33M0R_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module BEM2RA$func( OA1, OA2, Z, M0, M1, M2);
input M0, M1, M2;
output OA1, OA2, Z;

	BEM2RA_udp_0(OA1,M0,M1,M2); 

	BEM2RA_udp_1(OA2,M0,M1,M2); 

	ADHCM2R_udp_1(Z,M0,M1); 
endmodule
`endcelldefine
`celldefine
module BEM4RA$func( OA1, OA2, Z, M0, M1, M2);
input M0, M1, M2;
output OA1, OA2, Z;

	BEM2RA_udp_0(OA1,M0,M1,M2); 

	BEM2RA_udp_1(OA2,M0,M1,M2); 

	ADHCM2R_udp_1(Z,M0,M1); 
endmodule
`endcelldefine
`celldefine
module BEM8RA$func( OA1, OA2, Z, M0, M1, M2);
input M0, M1, M2;
output OA1, OA2, Z;

	BEM2RA_udp_0(OA1,M0,M1,M2); 

	BEM2RA_udp_1(OA2,M0,M1,M2); 

	ADHCM2R_udp_1(Z,M0,M1); 
endmodule
`endcelldefine
`celldefine
module BEMXBM2R$func( PB, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output PB;

	BEMXBM2R_udp_0(PB,M0,OA1,Z,OA2,M1); 
endmodule
`endcelldefine
`celldefine
module BEMXBM4R$func( PB, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output PB;

	BEMXBM2R_udp_0(PB,M0,OA1,Z,OA2,M1); 
endmodule
`endcelldefine
`celldefine
module BEMXM2RA$func( P, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output P;

	BEMXM2RA_udp_0(P,M0,OA1,Z,OA2,M1); 
endmodule
`endcelldefine
`celldefine
module BEMXM4RA$func( P, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output P;

	BEMXM2RA_udp_0(P,M0,OA1,Z,OA2,M1); 
endmodule
`endcelldefine
`celldefine
module BEMXM8RA$func( P, M0, M1, OA1, OA2, Z);
input M0, M1, OA1, OA2, Z;
output P;

	BEMXM2RA_udp_0(P,M0,OA1,Z,OA2,M1); 
endmodule
`endcelldefine
`celldefine
module BUFM10R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM12R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM14R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM16R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM18R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM20R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM22RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM24R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM26RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM2R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM32RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM3R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM40RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM48RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM4R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM5R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM6R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFM8R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module BUFTM0R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_1(MGM_WB_1,E);

	bufif0 MGM_BG_2(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM12R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM16R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM1R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM20R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM22RA$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM24RA$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM2R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM32RA$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM3R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM40RA$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM48RA$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM4R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM6R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module BUFTM8R$func( Z, A, E);
input A, E;
output Z;

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,A,E); 

	not MGM_BG_0(MGM_WB_1,E);

	bufif0 MGM_BG_1(Z,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module CKAN2M12R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKAN2M16RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKAN2M2R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKAN2M3R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKAN2M4R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKAN2M6R$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKAN2M8RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKBUFM12R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM16R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM1R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM20R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM22RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM24R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM26RA$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM2R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM32R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM3R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM40R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM48R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM4R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM6R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKBUFM8R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM12R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM16R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM1R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM20R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM22RA$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM24R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM26RA$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM2R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM32R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM3R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM40R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM48R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM4R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM6R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKINVM8R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module CKMUX2M12R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKMUX2M16RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKMUX2M2R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKMUX2M3R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKMUX2M4R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKMUX2M6R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKMUX2M8R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module CKND2M12R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKND2M16RA$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKND2M2R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKND2M4R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKND2M6RA$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKND2M8R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKXOR2M12RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKXOR2M1RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKXOR2M2RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKXOR2M4RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module CKXOR2M8RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module DEL1M1R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL1M4R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL2M1R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL2M4R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL3M1R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL3M4R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL4M1R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DEL4M4R$func( Z, A);
input A;
output Z;

	buf MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module DFAQM1RA$func( Q, A, B, CK,notifier);
input A, B, CK;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,A,B); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFAQM2RA$func( Q, A, B, CK,notifier);
input A, B, CK;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,A,B); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFAQM4RA$func( Q, A, B, CK,notifier);
input A, B, CK;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,A,B); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFAQM6RA$func( Q, A, B, CK,notifier);
input A, B, CK;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,A,B); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFAQM8RA$func( Q, A, B, CK,notifier);
input A, B, CK;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,A,B); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCM1RA$func( Q, QB, CKB, D,notifier);
input CKB, D;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCM2RA$func( Q, QB, CKB, D,notifier);
input CKB, D;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCM4RA$func( Q, QB, CKB, D,notifier);
input CKB, D;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCM8RA$func( Q, QB, CKB, D,notifier);
input CKB, D;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCQM1RA$func( Q, CKB, D,notifier);
input CKB, D;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQM2RA$func( Q, CKB, D,notifier);
input CKB, D;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQM4RA$func( Q, CKB, D,notifier);
input CKB, D;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQM8RA$func( Q, CKB, D,notifier);
input CKB, D;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRM1RA$func( Q, CKB, D, RB,notifier);
input CKB, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRM2RA$func( Q, CKB, D, RB,notifier);
input CKB, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRM4RA$func( Q, CKB, D, RB,notifier);
input CKB, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRM8RA$func( Q, CKB, D, RB,notifier);
input CKB, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRSM1RA$func( Q, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRSM2RA$func( Q, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRSM4RA$func( Q, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQRSM8RA$func( Q, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQSM1RA$func( Q, CKB, D, SB,notifier);
input CKB, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQSM2RA$func( Q, CKB, D, SB,notifier);
input CKB, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQSM4RA$func( Q, CKB, D, SB,notifier);
input CKB, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCQSM8RA$func( Q, CKB, D, SB,notifier);
input CKB, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFCRM1RA$func( Q, QB, CKB, D, RB,notifier);
input CKB, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRM2RA$func( Q, QB, CKB, D, RB,notifier);
input CKB, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRM4RA$func( Q, QB, CKB, D, RB,notifier);
input CKB, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRM8RA$func( Q, QB, CKB, D, RB,notifier);
input CKB, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRSM1RA$func( Q, QB, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRSM2RA$func( Q, QB, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRSM4RA$func( Q, QB, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCRSM8RA$func( Q, QB, CKB, D, RB, SB,notifier);
input CKB, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCSM1RA$func( Q, QB, CKB, D, SB,notifier);
input CKB, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCSM2RA$func( Q, QB, CKB, D, SB,notifier);
input CKB, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCSM4RA$func( Q, QB, CKB, D, SB,notifier);
input CKB, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFCSM8RA$func( Q, QB, CKB, D, SB,notifier);
input CKB, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEM1RA$func( Q, QB, CK, D, E,notifier);
input CK, D, E;
output Q, QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEM2RA$func( Q, QB, CK, D, E,notifier);
input CK, D, E;
output Q, QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEM4RA$func( Q, QB, CK, D, E,notifier);
input CK, D, E;
output Q, QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEM8RA$func( Q, QB, CK, D, E,notifier);
input CK, D, E;
output Q, QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEQBM1RA$func( QB, CK, D, E,notifier);
input CK, D, E;
output QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEQBM2RA$func( QB, CK, D, E,notifier);
input CK, D, E;
output QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEQBM4RA$func( QB, CK, D, E,notifier);
input CK, D, E;
output QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEQBM8RA$func( QB, CK, D, E,notifier);
input CK, D, E;
output QB;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEQM0RA$func( Q, CK, D, E,notifier);
input CK, D, E;
output Q;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQM1RA$func( Q, CK, D, E,notifier);
input CK, D, E;
output Q;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQM2RA$func( Q, CK, D, E,notifier);
input CK, D, E;
output Q;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQM4RA$func( Q, CK, D, E,notifier);
input CK, D, E;
output Q;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQM8RA$func( Q, CK, D, E,notifier);
input CK, D, E;
output Q;
input notifier;

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQRM1RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQRM2RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQRM4RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQRM8RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQZRM1RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQZRM2RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQZRM4RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFEQZRM8RA$func( Q, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFERM1RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFERM2RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFERM4RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFERM8RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	DFEM1RA_udp_0(MGM_D,D,E,IQ); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEZRM1RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEZRM2RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEZRM4RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFEZRM8RA$func( Q, QB, CK, D, E, RB,notifier);
input CK, D, E, RB;
output Q, QB;
input notifier;

	DFEQZRM1RA_udp_0(MGM_D,D,E,RB,IQ); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFM1RA$func( Q, QB, CK, D,notifier);
input CK, D;
output Q, QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFM2RA$func( Q, QB, CK, D,notifier);
input CK, D;
output Q, QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFM4RA$func( Q, QB, CK, D,notifier);
input CK, D;
output Q, QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFM8RA$func( Q, QB, CK, D,notifier);
input CK, D;
output Q, QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFMM1RA$func( Q, QB, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q, QB;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFMM2RA$func( Q, QB, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q, QB;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFMM4RA$func( Q, QB, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q, QB;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFMM8RA$func( Q, QB, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q, QB;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFMQM1RA$func( Q, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFMQM2RA$func( Q, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFMQM4RA$func( Q, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFMQM8RA$func( Q, CK, D1, D2, S,notifier);
input CK, D1, D2, S;
output Q;
input notifier;

	DFMM1RA_udp_0(MGM_D,D1,S,D2); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQBM1RA$func( QB, CK, D,notifier);
input CK, D;
output QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBM2RA$func( QB, CK, D,notifier);
input CK, D;
output QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBM4RA$func( QB, CK, D,notifier);
input CK, D;
output QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBM8RA$func( QB, CK, D,notifier);
input CK, D;
output QB;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBRM1RA$func( QB, CK, D, RB,notifier);
input CK, D, RB;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBRM2RA$func( QB, CK, D, RB,notifier);
input CK, D, RB;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBRM4RA$func( QB, CK, D, RB,notifier);
input CK, D, RB;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQBRM8RA$func( QB, CK, D, RB,notifier);
input CK, D, RB;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFQM1RA$func( Q, CK, D,notifier);
input CK, D;
output Q;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQM2RA$func( Q, CK, D,notifier);
input CK, D;
output Q;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQM4RA$func( Q, CK, D,notifier);
input CK, D;
output Q;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQM8RA$func( Q, CK, D,notifier);
input CK, D;
output Q;
input notifier;

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRM1RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRM2RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRM4RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRM8RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRSM1RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRSM2RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRSM4RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQRSM8RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQSM1RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQSM2RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQSM4RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQSM8RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRM1RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRM2RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRM4RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRM8RA$func( Q, CK, D, RB,notifier);
input CK, D, RB;
output Q;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRSM1RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRSM2RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRSM4RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZRSM8RA$func( Q, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZSM1RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZSM2RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZSM4RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFQZSM8RA$func( Q, CK, D, SB,notifier);
input CK, D, SB;
output Q;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module DFRM1RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRM2RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRM4RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRM8RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRSM1RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRSM2RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRSM4RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFRSM8RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFSM1RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFSM2RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFSM4RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFSM8RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRM1RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRM2RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRM4RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRM8RA$func( Q, QB, CK, D, RB,notifier);
input CK, D, RB;
output Q, QB;
input notifier;

	ADHM1RA_udp_0(MGM_D,D,RB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRSM1RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRSM2RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRSM4RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZRSM8RA$func( Q, QB, CK, D, RB, SB,notifier);
input CK, D, RB, SB;
output Q, QB;
input notifier;

	DFQZRSM1RA_udp_0(MGM_D,D,RB,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZSM1RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZSM2RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZSM4RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module DFZSM8RA$func( Q, QB, CK, D, SB,notifier);
input CK, D, SB;
output Q, QB;
input notifier;

	DFQZSM1RA_udp_0(MGM_D,D,SB); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module INVM0R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM10R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM12R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM14R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM16R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM18R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM1R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM20R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM22RA$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM24R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM26RA$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM2R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM32R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM3R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM40R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM48R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM4R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM5R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM6R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module INVM8R$func( Z, A);
input A;
output Z;

	not MGM_BG_0(Z,A);
endmodule
`endcelldefine
`celldefine
module LACM1RA$func( Q, QB, D, GB,notifier);
input D, GB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACM2RA$func( Q, QB, D, GB,notifier);
input D, GB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACM4RA$func( Q, QB, D, GB,notifier);
input D, GB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACM8RA$func( Q, QB, D, GB,notifier);
input D, GB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACQM1RA$func( Q, D, GB,notifier);
input D, GB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQM2RA$func( Q, D, GB,notifier);
input D, GB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQM4RA$func( Q, D, GB,notifier);
input D, GB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQM8RA$func( Q, D, GB,notifier);
input D, GB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRM1RA$func( Q, D, GB, RB,notifier);
input D, GB, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRM2RA$func( Q, D, GB, RB,notifier);
input D, GB, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRM4RA$func( Q, D, GB, RB,notifier);
input D, GB, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRM8RA$func( Q, D, GB, RB,notifier);
input D, GB, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRSM1RA$func( Q, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRSM2RA$func( Q, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRSM4RA$func( Q, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQRSM8RA$func( Q, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQSM1RA$func( Q, D, GB, SB,notifier);
input D, GB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQSM2RA$func( Q, D, GB, SB,notifier);
input D, GB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQSM4RA$func( Q, D, GB, SB,notifier);
input D, GB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACQSM8RA$func( Q, D, GB, SB,notifier);
input D, GB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LACRM1RA$func( Q, QB, D, GB, RB,notifier);
input D, GB, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRM2RA$func( Q, QB, D, GB, RB,notifier);
input D, GB, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRM4RA$func( Q, QB, D, GB, RB,notifier);
input D, GB, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRM8RA$func( Q, QB, D, GB, RB,notifier);
input D, GB, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRSM1RA$func( Q, QB, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRSM2RA$func( Q, QB, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRSM4RA$func( Q, QB, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACRSM8RA$func( Q, QB, D, GB, RB, SB,notifier);
input D, GB, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,MGM_EN,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACSM1RA$func( Q, QB, D, GB, SB,notifier);
input D, GB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACSM2RA$func( Q, QB, D, GB, SB,notifier);
input D, GB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACSM4RA$func( Q, QB, D, GB, SB,notifier);
input D, GB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LACSM8RA$func( Q, QB, D, GB, SB,notifier);
input D, GB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_EN,GB);

	not MGM_BG_1(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,MGM_EN,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,MGM_EN,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LAGCECSM12RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM12RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM16RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM16RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM24RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM24RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM2RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM2RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM32RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM32RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM40RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM40RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM48RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM48RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM4RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM4RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM6RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM6RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCECSM8RA$func( GCK, CKB, E, SE,notifier);
input CKB, E, SE;
output GCK;
input notifier;

	LAGCECSM8RA_statetable_ENL(ENL,CKB,E,SE);
	DFQZSM1RA_udp_0(GCK,CKB,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM12R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM12R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM16R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM16R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM20R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM20R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM2R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM2R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM3R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM3R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM4R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM4R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM6R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM6R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEM8R$func( GCK, CK, E,notifier);
input CK, E;
output GCK;
input notifier;

	LAGCEM8R_statetable_ENL(ENL,CK,E);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM12R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM12R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM16R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM16R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM20R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM20R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM2R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM2R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM3R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM3R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM4R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM4R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM6R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM6R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPM8R$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCEPM8R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 
endmodule
`endcelldefine
`celldefine
module LAGCEPOM12R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM12R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM16R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM16R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM20R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM20R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM2R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM2R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM3R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM3R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM4R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM4R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM6R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM6R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCEPOM8R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCEPOM8R_statetable_ENL(ENL,CK,E);
	LAGCEPM12R_udp_0(GCK,CK,ENL,SE); 

	buf MGM_BG_0(OBS,ENL);
endmodule
`endcelldefine
`celldefine
module LAGCESM12RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM12RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM16RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM16RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM24RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM24RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM2RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM2RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM32RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM32RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM40RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM40RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM48RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM48RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM4RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM4RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM6RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM6RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESM8RA$func( GCK, CK, E, SE,notifier);
input CK, E, SE;
output GCK;
input notifier;

	LAGCESM8RA_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 
endmodule
`endcelldefine
`celldefine
module LAGCESOM12R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM12R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM16R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM16R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM20R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM20R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM2R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM2R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM3R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM3R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM4R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM4R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM6R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM6R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAGCESOM8R$func( GCK, OBS, CK, E, SE,notifier);
input CK, E, SE;
output GCK, OBS;
input notifier;

	LAGCESOM8R_statetable_ENL(ENL,CK,E,SE);
	ADHM1RA_udp_0(GCK,CK,ENL); 

	buf MGM_BG_0(OBS,E);
endmodule
`endcelldefine
`celldefine
module LAM1RA$func( Q, QB, D, G,notifier);
input D, G;
output Q, QB;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LAM2RA$func( Q, QB, D, G,notifier);
input D, G;
output Q, QB;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LAM4RA$func( Q, QB, D, G,notifier);
input D, G;
output Q, QB;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LAM8RA$func( Q, QB, D, G,notifier);
input D, G;
output Q, QB;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LAQM1RA$func( Q, D, G,notifier);
input D, G;
output Q;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQM2RA$func( Q, D, G,notifier);
input D, G;
output Q;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQM4RA$func( Q, D, G,notifier);
input D, G;
output Q;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQM8RA$func( Q, D, G,notifier);
input D, G;
output Q;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,G,D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRM1RA$func( Q, D, G, RB,notifier);
input D, G, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRM2RA$func( Q, D, G, RB,notifier);
input D, G, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRM4RA$func( Q, D, G, RB,notifier);
input D, G, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRM8RA$func( Q, D, G, RB,notifier);
input D, G, RB;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRSM1RA$func( Q, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRSM2RA$func( Q, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRSM4RA$func( Q, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQRSM8RA$func( Q, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQSM1RA$func( Q, D, G, SB,notifier);
input D, G, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQSM2RA$func( Q, D, G, SB,notifier);
input D, G, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQSM4RA$func( Q, D, G, SB,notifier);
input D, G, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LAQSM8RA$func( Q, D, G, SB,notifier);
input D, G, SB;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module LARM1RA$func( Q, QB, D, G, RB,notifier);
input D, G, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARM2RA$func( Q, QB, D, G, RB,notifier);
input D, G, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARM4RA$func( Q, QB, D, G, RB,notifier);
input D, G, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARM8RA$func( Q, QB, D, G, RB,notifier);
input D, G, RB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	MGM_IQ_LATCH_UDP(IQ,MGM_C,1'b0,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,MGM_C,1'b0,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARSM1RA$func( Q, QB, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARSM2RA$func( Q, QB, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARSM4RA$func( Q, QB, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LARSM8RA$func( Q, QB, D, G, RB, SB,notifier);
input D, G, RB, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	MGM_H_IQ_LATCH_UDP(IQ,MGM_C,MGM_P,G,D,notifier);

	MGM_L_IQN_LATCH_UDP(IQN,MGM_C,MGM_P,G,D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LASM1RA$func( Q, QB, D, G, SB,notifier);
input D, G, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LASM2RA$func( Q, QB, D, G, SB,notifier);
input D, G, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LASM4RA$func( Q, QB, D, G, SB,notifier);
input D, G, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module LASM8RA$func( Q, QB, D, G, SB,notifier);
input D, G, SB;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	MGM_IQ_LATCH_UDP(IQ,1'b0,MGM_P,G,D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,MGM_P,G,D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module MAO222M1RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AD42M2RA_udp_1(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAO222M2RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AD42M2RA_udp_1(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAO222M4RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AD42M2RA_udp_1(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAO222M8RA$func( Z, A, B, C);
input A, B, C;
output Z;

	AD42M2RA_udp_1(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAOI2223M1RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	MAOI2223M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MAOI2223M2RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	MAOI2223M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MAOI2223M4RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	MAOI2223M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MAOI2223M8RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	MAOI2223M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MAOI222M1RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADCSOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAOI222M2RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADCSOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAOI222M4RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADCSOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAOI222M8RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADCSOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module MAOI22M1RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22B20M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module MAOI22M2RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22B20M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module MAOI22M4RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22B20M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module MAOI22M8RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	AOI22B20M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module MOAI22M1RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	MOAI22M1RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module MOAI22M2RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	MOAI22M1RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module MOAI22M4RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	MOAI22M1RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module MOAI22M8RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	MOAI22M1RA_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module MUX2M0RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M12RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M1RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M2RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M3RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M4RA$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M6R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX2M8R$func( Z, A, B, S);
input A, B, S;
output Z;

	CKMUX2M12R_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MUX3M0RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MUX3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MUX3M1RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MUX3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MUX3M2RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MUX3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MUX3M4RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MUX3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MUX3M8RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MUX3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MUX4M0RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MUX4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MUX4M1RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MUX4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MUX4M2RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MUX4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MUX4M4R$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MUX4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MUX4M8RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MUX4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MXB2M0RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB2M1RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB2M2RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB2M3RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB2M4RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB2M6RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB2M8RA$func( Z, A, B, S);
input A, B, S;
output Z;

	MXB2M0RA_udp_0(Z,A,S,B); 
endmodule
`endcelldefine
`celldefine
module MXB3M0RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MXB3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MXB3M1RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MXB3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MXB3M2RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MXB3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MXB3M4RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MXB3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MXB3M8RA$func( Z, A, B, C, S0, S1);
input A, B, C, S0, S1;
output Z;

	MXB3M0RA_udp_0(Z,A,S0,S1,B,C); 
endmodule
`endcelldefine
`celldefine
module MXB4M0RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MXB4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MXB4M1RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MXB4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MXB4M2RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MXB4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MXB4M4RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MXB4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MXB4M6RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MXB4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module MXB4M8RA$func( Z, A, B, C, D, S0, S1);
input A, B, C, D, S0, S1;
output Z;

	MXB4M0RA_udp_0(Z,A,S0,S1,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND2B1M0R$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M12RA$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M16RA$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M1R$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M2R$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M4R$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M6RA$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2B1M8R$func( Z, B, NA);
input B, NA;
output Z;

	ND2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module ND2M0R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M12RA$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M16RA$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M1R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M2R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M3R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M4R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M5R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M6R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND2M8R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module ND3B1M0R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3B1M12RA$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3B1M1R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3B1M2R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3B1M4R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3B1M6RA$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3B1M8RA$func( Z, B, C, NA);
input B, C, NA;
output Z;

	ND3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module ND3M0R$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M12RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M16RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M1R$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M2R$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M3R$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M4RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M6RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND3M8RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ND3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module ND4B1M0R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	ND4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module ND4B1M1R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	ND4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module ND4B1M2R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	ND4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module ND4B1M4R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	ND4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module ND4B1M6RA$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	ND4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module ND4B1M8RA$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	ND4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module ND4B2M0R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	ND4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module ND4B2M1R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	ND4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module ND4B2M2R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	ND4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module ND4B2M4R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	ND4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module ND4B2M8RA$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	ND4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module ND4M0R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND4M16RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND4M1R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND4M2R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND4M4R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND4M6R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module ND4M8R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	ND4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR2B1M0R$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M12RA$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M16RA$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M1R$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M2R$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M4R$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M6RA$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2B1M8R$func( Z, B, NA);
input B, NA;
output Z;

	NR2B1M0R_udp_0(Z,B,NA); 
endmodule
`endcelldefine
`celldefine
module NR2M0R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M12RA$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M16RA$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M1R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M2R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M3R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M4R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M5R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M6R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR2M8R$func( Z, A, B);
input A, B;
output Z;

	ADCSIOM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module NR3B1M0R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	NR3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module NR3B1M1R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	NR3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module NR3B1M2R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	NR3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module NR3B1M4R$func( Z, B, C, NA);
input B, C, NA;
output Z;

	NR3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module NR3B1M8RA$func( Z, B, C, NA);
input B, C, NA;
output Z;

	NR3B1M0R_udp_0(Z,B,C,NA); 
endmodule
`endcelldefine
`celldefine
module NR3M0R$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR3M16RA$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR3M1R$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR3M2R$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR3M4R$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR3M6R$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR3M8R$func( Z, A, B, C);
input A, B, C;
output Z;

	NR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module NR4B1M0R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	NR4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module NR4B1M1R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	NR4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module NR4B1M2R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	NR4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module NR4B1M4R$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	NR4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module NR4B1M8RA$func( Z, B, C, D, NA);
input B, C, D, NA;
output Z;

	NR4B1M0R_udp_0(Z,B,C,D,NA); 
endmodule
`endcelldefine
`celldefine
module NR4B2M0R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	NR4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module NR4B2M1R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	NR4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module NR4B2M2R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	NR4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module NR4B2M4R$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	NR4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module NR4B2M8RA$func( Z, C, D, NA, NB);
input C, D, NA, NB;
output Z;

	NR4B2M0R_udp_0(Z,C,D,NA,NB); 
endmodule
`endcelldefine
`celldefine
module NR4M0R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR4M16RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR4M1R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR4M2R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR4M4RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR4M6R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module NR4M8RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	NR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OA211M12RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OA211M12RA_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module OA211M1RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OA211M12RA_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module OA211M2RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OA211M12RA_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module OA211M4RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OA211M12RA_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module OA211M6RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OA211M12RA_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module OA211M8RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OA211M12RA_udp_0(Z,A1,B,C,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M0RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M12RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M16RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M1RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M2RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M4RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M6RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA21M8RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OA21M0RA_udp_0(Z,A1,B,A2); 
endmodule
`endcelldefine
`celldefine
module OA221M1RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OA221M1RA_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA221M2RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OA221M1RA_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA221M4RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OA221M1RA_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA221M8RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OA221M1RA_udp_0(Z,A1,B1,C,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA222M1RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OA222M1RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA222M2RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OA222M1RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA222M4RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OA222M1RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA222M8RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OA222M1RA_udp_0(Z,A1,B1,C1,C2,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M0R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M12RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M16RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M1R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M2R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M4R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M6RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA22M8RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OA22M0R_udp_0(Z,A1,B1,B2,A2); 
endmodule
`endcelldefine
`celldefine
module OA31M1RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OA31M1RA_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA31M2RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OA31M1RA_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA31M4RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OA31M1RA_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA31M8RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OA31M1RA_udp_0(Z,A1,B,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA32M1RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OA32M1RA_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA32M2RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OA32M1RA_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA32M4RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OA32M1RA_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA32M8RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OA32M1RA_udp_0(Z,A1,B1,B2,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA33M1RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OA33M1RA_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA33M2RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OA33M1RA_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA33M4RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OA33M1RA_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OA33M8RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OA33M1RA_udp_0(Z,A1,B1,B2,B3,A2,A3); 
endmodule
`endcelldefine
`celldefine
module OAI211B100M0R$func( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

	OAI211B100M0R_udp_0(Z,A1,NA2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211B100M1R$func( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

	OAI211B100M0R_udp_0(Z,A1,NA2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211B100M2R$func( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

	OAI211B100M0R_udp_0(Z,A1,NA2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211B100M4R$func( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

	OAI211B100M0R_udp_0(Z,A1,NA2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211B100M8RA$func( Z, A1, B, C, NA2);
input A1, B, C, NA2;
output Z;

	OAI211B100M0R_udp_0(Z,A1,NA2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211M0R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OAI211M0R_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211M1R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OAI211M0R_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211M2R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OAI211M0R_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211M4R$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OAI211M0R_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211M6RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OAI211M0R_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI211M8RA$func( Z, A1, A2, B, C);
input A1, A2, B, C;
output Z;

	OAI211M0R_udp_0(Z,A1,A2,B,C); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M0R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M12RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M16RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M1R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M2R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M4R$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M6RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B01M8RA$func( Z, A1, A2, NB);
input A1, A2, NB;
output Z;

	BEM2RA_udp_1(Z,A1,A2,NB); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M0R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M12RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M16RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M1R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M2R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M4R$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M6RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B10M8RA$func( Z, A1, B, NA2);
input A1, B, NA2;
output Z;

	OAI21B10M0R_udp_0(Z,A1,NA2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M0R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M12RA$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M1R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M2R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M4R$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M6RA$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21B20M8RA$func( Z, B, NA1, NA2);
input B, NA1, NA2;
output Z;

	OAI21B20M0R_udp_0(Z,B,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI21M0R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M12RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M16RA$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M1R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M2R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M3R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M4R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M6R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI21M8R$func( Z, A1, A2, B);
input A1, A2, B;
output Z;

	OAI21M0R_udp_0(Z,A1,A2,B); 
endmodule
`endcelldefine
`celldefine
module OAI221M0R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OAI221M0R_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module OAI221M1R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OAI221M0R_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module OAI221M2R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OAI221M0R_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module OAI221M4R$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OAI221M0R_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module OAI221M6RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OAI221M0R_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module OAI221M8RA$func( Z, A1, A2, B1, B2, C);
input A1, A2, B1, B2, C;
output Z;

	OAI221M0R_udp_0(Z,A1,A2,B1,B2,C); 
endmodule
`endcelldefine
`celldefine
module OAI222M0RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OAI222M0RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module OAI222M1RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OAI222M0RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module OAI222M2RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OAI222M0RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module OAI222M4R$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OAI222M0RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module OAI222M6RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OAI222M0RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module OAI222M8RA$func( Z, A1, A2, B1, B2, C1, C2);
input A1, A2, B1, B2, C1, C2;
output Z;

	OAI222M0RA_udp_0(Z,A1,A2,B1,B2,C1,C2); 
endmodule
`endcelldefine
`celldefine
module OAI22B10M0R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	OAI22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22B10M1R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	OAI22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22B10M2R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	OAI22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22B10M4R$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	OAI22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22B10M8RA$func( Z, A1, B1, B2, NA2);
input A1, B1, B2, NA2;
output Z;

	OAI22B10M0R_udp_0(Z,A1,NA2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22B20M0R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	MOAI22M1RA_udp_0(Z,B1,B2,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI22B20M1R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	MOAI22M1RA_udp_0(Z,B1,B2,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI22B20M2R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	MOAI22M1RA_udp_0(Z,B1,B2,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI22B20M4R$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	MOAI22M1RA_udp_0(Z,B1,B2,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI22B20M8RA$func( Z, B1, B2, NA1, NA2);
input B1, B2, NA1, NA2;
output Z;

	MOAI22M1RA_udp_0(Z,B1,B2,NA1,NA2); 
endmodule
`endcelldefine
`celldefine
module OAI22M0R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M12RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M16RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M1R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M2R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M4R$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M6RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI22M8RA$func( Z, A1, A2, B1, B2);
input A1, A2, B1, B2;
output Z;

	OAI22M0R_udp_0(Z,A1,A2,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI31M0R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OAI31M0R_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module OAI31M1R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OAI31M0R_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module OAI31M2R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OAI31M0R_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module OAI31M4R$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OAI31M0R_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module OAI31M8RA$func( Z, A1, A2, A3, B);
input A1, A2, A3, B;
output Z;

	OAI31M0R_udp_0(Z,A1,A2,A3,B); 
endmodule
`endcelldefine
`celldefine
module OAI32M0R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OAI32M0R_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI32M1R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OAI32M0R_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI32M2R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OAI32M0R_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI32M4R$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OAI32M0R_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI32M8RA$func( Z, A1, A2, A3, B1, B2);
input A1, A2, A3, B1, B2;
output Z;

	OAI32M0R_udp_0(Z,A1,A2,A3,B1,B2); 
endmodule
`endcelldefine
`celldefine
module OAI33M0R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OAI33M0R_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module OAI33M1R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OAI33M0R_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module OAI33M2R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OAI33M0R_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module OAI33M4R$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OAI33M0R_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module OAI33M8RA$func( Z, A1, A2, A3, B1, B2, B3);
input A1, A2, A3, B1, B2, B3;
output Z;

	OAI33M0R_udp_0(Z,A1,A2,A3,B1,B2,B3); 
endmodule
`endcelldefine
`celldefine
module OR2M0R$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M12RA$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M16RA$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M1R$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M22RA$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M2R$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M4R$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M6R$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR2M8R$func( Z, A, B);
input A, B;
output Z;

	OR2M0R_udp_0(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module OR3M0R$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M12RA$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M16RA$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M1R$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M2R$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M4R$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M6R$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR3M8RA$func( Z, A, B, C);
input A, B, C;
output Z;

	OR3M0R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module OR4M0R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M12RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M16RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M1R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M2R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M4RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M6R$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR4M8RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	OR4M0R_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module OR6M12RA$func( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

	OR6M12RA_udp_0(Z,A,B,C,D,E,F); 
endmodule
`endcelldefine
`celldefine
module OR6M1RA$func( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

	OR6M12RA_udp_0(Z,A,B,C,D,E,F); 
endmodule
`endcelldefine
`celldefine
module OR6M2RA$func( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

	OR6M12RA_udp_0(Z,A,B,C,D,E,F); 
endmodule
`endcelldefine
`celldefine
module OR6M4RA$func( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

	OR6M12RA_udp_0(Z,A,B,C,D,E,F); 
endmodule
`endcelldefine
`celldefine
module OR6M6RA$func( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

	OR6M12RA_udp_0(Z,A,B,C,D,E,F); 
endmodule
`endcelldefine
`celldefine
module OR6M8RA$func( Z, A, B, C, D, E, F);
input A, B, C, D, E, F;
output Z;

	OR6M12RA_udp_0(Z,A,B,C,D,E,F); 
endmodule
`endcelldefine
`celldefine
module REG1M1R$func( RQB, RD, RG, RGB, WE,notifier);
input RD, RG, RGB, WE;
output RQB;
input notifier;

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,WE,RD,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,WE,RD,notifier);

	wire MGM_WB_0;

	wire MGM_WB_1;

	REG1M1R_udp_0(MGM_WB_0,IQN,RG,RGB); 

	ND2B1M0R_udp_0(MGM_WB_1,RG,RGB); 

	bufif0 MGM_BG_1(RQB,MGM_WB_0,MGM_WB_1);
endmodule
`endcelldefine
`celldefine
module REG2M1R$func( RQ1B, RQ2B, RD, RG1, RG2, WE,notifier);
input RD, RG1, RG2, WE;
output RQ1B, RQ2B;
input notifier;

	not MGM_BG_0(MGM_D,RD);

	MGM_IQ_LATCH_UDP(IQ,1'b0,1'b0,WE,MGM_D,notifier);

	MGM_IQN_LATCH_UDP(IQN,1'b0,1'b0,WE,MGM_D,notifier);

	wire MGM_WB_0;

	wire MGM_WB_1;

	BUFTM0R_udp_0(MGM_WB_0,IQ,RG1); 

	not MGM_BG_1(MGM_WB_1,RG1);

	bufif0 MGM_BG_2(RQ1B,MGM_WB_0,MGM_WB_1);

	wire MGM_WB_2;

	wire MGM_WB_3;

	BUFTM0R_udp_0(MGM_WB_2,IQ,RG2); 

	not MGM_BG_3(MGM_WB_3,RG2);

	bufif0 MGM_BG_4(RQ2B,MGM_WB_2,MGM_WB_3);
endmodule
`endcelldefine
`celldefine
module REGKM1R$func( RQB, RD);
input RD;
output RQB;

	not MGM_BG_0(RQB,RD);
endmodule
`endcelldefine
`celldefine
module REGKM2R$func( RQB, RD);
input RD;
output RQB;

	not MGM_BG_0(RQB,RD);
endmodule
`endcelldefine
`celldefine
module REGKM4R$func( RQB, RD);
input RD;
output RQB;

	not MGM_BG_0(RQB,RD);
endmodule
`endcelldefine
`celldefine
module SDFAQM1RA$func( Q, A, B, CK, SD, SE,notifier);
input A, B, CK, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,A,B,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFAQM2RA$func( Q, A, B, CK, SD, SE,notifier);
input A, B, CK, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,A,B,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFAQM4RA$func( Q, A, B, CK, SD, SE,notifier);
input A, B, CK, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,A,B,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFAQM6RA$func( Q, A, B, CK, SD, SE,notifier);
input A, B, CK, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,A,B,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFAQM8RA$func( Q, A, B, CK, SD, SE,notifier);
input A, B, CK, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,A,B,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCM1RA$func( Q, QB, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCM2RA$func( Q, QB, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCM4RA$func( Q, QB, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCM8RA$func( Q, QB, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCQM1RA$func( Q, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQM2RA$func( Q, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQM4RA$func( Q, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQM8RA$func( Q, CKB, D, SD, SE,notifier);
input CKB, D, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRM1RA$func( Q, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRM2RA$func( Q, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRM4RA$func( Q, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRM8RA$func( Q, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRSM1RA$func( Q, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRSM2RA$func( Q, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRSM4RA$func( Q, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQRSM8RA$func( Q, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQSM1RA$func( Q, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQSM2RA$func( Q, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQSM4RA$func( Q, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCQSM8RA$func( Q, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFCRM1RA$func( Q, QB, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRM2RA$func( Q, QB, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRM4RA$func( Q, QB, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRM8RA$func( Q, QB, CKB, D, RB, SD, SE,notifier);
input CKB, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRSM1RA$func( Q, QB, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRSM2RA$func( Q, QB, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRSM4RA$func( Q, QB, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCRSM8RA$func( Q, QB, CKB, D, RB, SB, SD, SE,notifier);
input CKB, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	not MGM_BG_2(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_3(Q,IQ);

	buf MGM_BG_4(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCSM1RA$func( Q, QB, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCSM2RA$func( Q, QB, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCSM4RA$func( Q, QB, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFCSM8RA$func( Q, QB, CKB, D, SB, SD, SE,notifier);
input CKB, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_CLK,CKB);

	not MGM_BG_1(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,MGM_CLK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEM1RA$func( Q, QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q, QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEM2RA$func( Q, QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q, QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEM4RA$func( Q, QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q, QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEM8RA$func( Q, QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q, QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEQBM1RA$func( QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEQBM2RA$func( QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEQBM4RA$func( QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEQBM8RA$func( QB, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output QB;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEQM0RA$func( Q, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQM1RA$func( Q, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQM2RA$func( Q, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQM4RA$func( Q, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQM8RA$func( Q, CK, D, E, SD, SE,notifier);
input CK, D, E, SD, SE;
output Q;
input notifier;

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQRM1RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQRM2RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQRM4RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQRM8RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQZRM1RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQZRM2RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQZRM4RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFEQZRM8RA$func( Q, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFERM1RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFERM2RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFERM4RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFERM8RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	SDFEM1RA_udp_0(MGM_D,D,E,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEZRM1RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEZRM2RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEZRM4RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFEZRM8RA$func( Q, QB, CK, D, E, RB, SD, SE,notifier);
input CK, D, E, RB, SD, SE;
output Q, QB;
input notifier;

	SDFEQZRM1RA_udp_0(MGM_D,D,E,RB,SE,IQ,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFM1RA$func( Q, QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q, QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFM2RA$func( Q, QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q, QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFM4RA$func( Q, QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q, QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFM8RA$func( Q, QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q, QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFMM1RA$func( Q, QB, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFMM2RA$func( Q, QB, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFMM4RA$func( Q, QB, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFMM8RA$func( Q, QB, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q, QB;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFMQM1RA$func( Q, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFMQM2RA$func( Q, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFMQM4RA$func( Q, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFMQM8RA$func( Q, CK, D1, D2, S, SD, SE,notifier);
input CK, D1, D2, S, SD, SE;
output Q;
input notifier;

	SDFMM1RA_udp_0(MGM_D,D1,S,SE,D2,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQBM1RA$func( QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBM2RA$func( QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBM4RA$func( QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBM8RA$func( QB, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output QB;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBRM1RA$func( QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBRM2RA$func( QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBRM4RA$func( QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQBRM8RA$func( QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFQM1RA$func( Q, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQM2RA$func( Q, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQM4RA$func( Q, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQM8RA$func( Q, CK, D, SD, SE,notifier);
input CK, D, SD, SE;
output Q;
input notifier;

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRM1RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRM2RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRM4RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRM8RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRSM1RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRSM2RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRSM4RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQRSM8RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_H_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQSM1RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQSM2RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQSM4RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQSM8RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRM1RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRM2RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRM4RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRM8RA$func( Q, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRSM1RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRSM2RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRSM4RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZRSM8RA$func( Q, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZSM1RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZSM2RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZSM4RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFQZSM8RA$func( Q, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);
endmodule
`endcelldefine
`celldefine
module SDFRM1RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRM2RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRM4RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRM8RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,MGM_C,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,MGM_C,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRSM1RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRSM2RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRSM4RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFRSM8RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	not MGM_BG_1(MGM_C,RB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_L_IQ_FF_UDP(IQ,MGM_C,MGM_P,CK,MGM_D,notifier);

	MGM_L_IQN_FF_UDP(IQN,MGM_C,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_2(Q,IQ);

	buf MGM_BG_3(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFSM1RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFSM2RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFSM4RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFSM8RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	not MGM_BG_0(MGM_P,SB);

	CKMUX2M12R_udp_0(MGM_D,D,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,MGM_P,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,MGM_P,CK,MGM_D,notifier);

	buf MGM_BG_1(Q,IQ);

	buf MGM_BG_2(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRM1RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRM2RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRM4RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRM8RA$func( Q, QB, CK, D, RB, SD, SE,notifier);
input CK, D, RB, SD, SE;
output Q, QB;
input notifier;

	SDFAQM1RA_udp_0(MGM_D,D,RB,SE,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRSM1RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRSM2RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRSM4RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZRSM8RA$func( Q, QB, CK, D, RB, SB, SD, SE,notifier);
input CK, D, RB, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZRSM1RA_udp_0(MGM_D,D,RB,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZSM1RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZSM2RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZSM4RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module SDFZSM8RA$func( Q, QB, CK, D, SB, SD, SE,notifier);
input CK, D, SB, SD, SE;
output Q, QB;
input notifier;

	SDFQZSM1RA_udp_0(MGM_D,D,SE,SB,SD); 

	MGM_IQ_FF_UDP(IQ,1'b0,1'b0,CK,MGM_D,notifier);

	MGM_IQN_FF_UDP(IQN,1'b0,1'b0,CK,MGM_D,notifier);

	buf MGM_BG_0(Q,IQ);

	buf MGM_BG_1(QB,IQN);
endmodule
`endcelldefine
`celldefine
module TIE0R$func( Z);
output Z;

	assign Z = 1'b0;
endmodule
`endcelldefine
`celldefine
module TIE1R$func( Z);
output Z;

	assign Z = 1'b1;
endmodule
`endcelldefine
`celldefine
module XNR2M0RA$func( Z, A, B);
input A, B;
output Z;

	ADHCM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XNR2M1RA$func( Z, A, B);
input A, B;
output Z;

	ADHCM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XNR2M2RA$func( Z, A, B);
input A, B;
output Z;

	ADHCM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XNR2M4RA$func( Z, A, B);
input A, B;
output Z;

	ADHCM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XNR2M6RA$func( Z, A, B);
input A, B;
output Z;

	ADHCM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XNR2M8RA$func( Z, A, B);
input A, B;
output Z;

	ADHCM2R_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XNR3M0RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCM2RA_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XNR3M1R$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCM2RA_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XNR3M2R$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCM2RA_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XNR3M4R$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCM2RA_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XNR3M6RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCM2RA_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XNR3M8RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCM2RA_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XNR4M1RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XNR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XNR4M2RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XNR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XNR4M4RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XNR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XNR4M8RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XNR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XOR2M0RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR2M1RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR2M2RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR2M3RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR2M4RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR2M6RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR2M8RA$func( Z, A, B);
input A, B;
output Z;

	ADHM1RA_udp_1(Z,A,B); 
endmodule
`endcelldefine
`celldefine
module XOR3M0RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCSIOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XOR3M1RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCSIOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XOR3M2RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCSIOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XOR3M4RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCSIOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XOR3M6RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCSIOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XOR3M8RA$func( Z, A, B, C);
input A, B, C;
output Z;

	ADFCSIOM2R_udp_0(Z,A,B,C); 
endmodule
`endcelldefine
`celldefine
module XOR4M1RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XOR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XOR4M2RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XOR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XOR4M4RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XOR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine
`celldefine
module XOR4M8RA$func( Z, A, B, C, D);
input A, B, C, D;
output Z;

	XOR4M1RA_udp_0(Z,A,B,C,D); 
endmodule
`endcelldefine

primitive AD42M2RA_udp_0(CO,A, B, C, D, ICI);
  output CO;
  input A, B, C, D, ICI;
  table
  //A, B, C, D, ICI: CO
    1  1  1  1  ?: 1;
    1  1  1  ?  1: 1;
    1  0  0  1  ?: 1;
    1  0  0  ?  1: 1;
    0  1  0  1  ?: 1;
    0  1  0  ?  1: 1;
    0  0  1  1  ?: 1;
    0  0  1  ?  1: 1;
    ?  ?  ?  1  1: 1;
    1  1  0  0  ?: 0;
    1  1  0  ?  0: 0;
    1  0  1  0  ?: 0;
    1  0  1  ?  0: 0;
    0  1  1  0  ?: 0;
    0  1  1  ?  0: 0;
    0  0  0  0  ?: 0;
    0  0  0  ?  0: 0;
    ?  ?  ?  0  0: 0;
  endtable
endprimitive

primitive AD42M2RA_udp_1(ICO,A, B, C);
  output ICO;
  input A, B, C;
  table
  //A, B, C: ICO
    1  1  ?: 1;
    1  ?  1: 1;
    ?  1  1: 1;
    0  0  ?: 0;
    0  ?  0: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive AD42M2RA_udp_2(S,A, B, C, D, ICI);
  output S;
  input A, B, C, D, ICI;
  table
  //A, B, C, D, ICI: S
    1  1  1  1  1: 1;
    1  1  1  0  0: 1;
    1  1  0  1  0: 1;
    1  1  0  0  1: 1;
    1  0  1  1  0: 1;
    1  0  1  0  1: 1;
    1  0  0  1  1: 1;
    1  0  0  0  0: 1;
    0  1  1  1  0: 1;
    0  1  1  0  1: 1;
    0  1  0  1  1: 1;
    0  1  0  0  0: 1;
    0  0  1  1  1: 1;
    0  0  1  0  0: 1;
    0  0  0  1  0: 1;
    0  0  0  0  1: 1;
    1  1  1  1  0: 0;
    1  1  1  0  1: 0;
    1  1  0  1  1: 0;
    1  1  0  0  0: 0;
    1  0  1  1  1: 0;
    1  0  1  0  0: 0;
    1  0  0  1  0: 0;
    1  0  0  0  1: 0;
    0  1  1  1  1: 0;
    0  1  1  0  0: 0;
    0  1  0  1  0: 0;
    0  1  0  0  1: 0;
    0  0  1  1  0: 0;
    0  0  1  0  1: 0;
    0  0  0  1  1: 0;
    0  0  0  0  0: 0;
  endtable
endprimitive

primitive ADCSCM2R_udp_0(CO0,A, B, NCI0);
  output CO0;
  input A, B, NCI0;
  table
  //A, B, NCI0: CO0
    1  1  ?: 1;
    1  ?  0: 1;
    ?  1  0: 1;
    0  0  ?: 0;
    0  ?  1: 0;
    ?  0  1: 0;
  endtable
endprimitive

primitive ADCSIOM2R_udp_0(CO0B,A, B);
  output CO0B;
  input A, B;
  table
  //A, B: CO0B
    0  ?: 1;
    ?  0: 1;
    1  1: 0;
  endtable
endprimitive

primitive ADCSIOM2R_udp_1(CO1B,A, B);
  output CO1B;
  input A, B;
  table
  //A, B: CO1B
    0  0: 1;
    1  ?: 0;
    ?  1: 0;
  endtable
endprimitive

primitive ADCSOM2R_udp_0(CO0B,A, B, CI0);
  output CO0B;
  input A, B, CI0;
  table
  //A, B, CI0: CO0B
    0  0  ?: 1;
    0  ?  0: 1;
    ?  0  0: 1;
    1  1  ?: 0;
    1  ?  1: 0;
    ?  1  1: 0;
  endtable
endprimitive

primitive ADFCM2RA_udp_0(S,A, B, NCI);
  output S;
  input A, B, NCI;
  table
  //A, B, NCI: S
    1  1  0: 1;
    1  0  1: 1;
    0  1  1: 1;
    0  0  0: 1;
    1  1  1: 0;
    1  0  0: 0;
    0  1  0: 0;
    0  0  1: 0;
  endtable
endprimitive

primitive ADFCSCM2RA_udp_0(S,A, B, CS, NCI1, NCI0);
  output S;
  input A, B, CS, NCI1, NCI0;
  table
  //A, B, CS, NCI1, NCI0: S
    1  1  1  0  ?: 1;
    1  1  0  ?  0: 1;
    1  1  ?  0  0: 1;
    1  0  1  1  ?: 1;
    1  0  0  ?  1: 1;
    1  0  ?  1  1: 1;
    0  1  1  1  ?: 1;
    0  1  0  ?  1: 1;
    0  1  ?  1  1: 1;
    0  0  1  0  ?: 1;
    0  0  0  ?  0: 1;
    0  0  ?  0  0: 1;
    1  1  1  1  ?: 0;
    1  1  0  ?  1: 0;
    1  1  ?  1  1: 0;
    1  0  1  0  ?: 0;
    1  0  0  ?  0: 0;
    1  0  ?  0  0: 0;
    0  1  1  0  ?: 0;
    0  1  0  ?  0: 0;
    0  1  ?  0  0: 0;
    0  0  1  1  ?: 0;
    0  0  0  ?  1: 0;
    0  0  ?  1  1: 0;
  endtable
endprimitive

primitive ADFCSIOM2R_udp_0(S,A, B, CS);
  output S;
  input A, B, CS;
  table
  //A, B, CS: S
    1  1  1: 1;
    1  0  0: 1;
    0  1  0: 1;
    0  0  1: 1;
    1  1  0: 0;
    1  0  1: 0;
    0  1  1: 0;
    0  0  0: 0;
  endtable
endprimitive

primitive ADFCSOM2RA_udp_0(S,A, B, CI0, CS, CI1);
  output S;
  input A, B, CI0, CS, CI1;
  table
  //A, B, CI0, CS, CI1: S
    1  1  1  0  ?: 1;
    1  1  ?  1  1: 1;
    1  0  0  0  ?: 1;
    1  0  ?  1  0: 1;
    0  1  0  0  ?: 1;
    0  1  ?  1  0: 1;
    0  0  1  0  ?: 1;
    0  0  ?  1  1: 1;
    1  1  0  0  ?: 0;
    1  1  ?  1  0: 0;
    1  0  1  0  ?: 0;
    1  0  ?  1  1: 0;
    0  1  1  0  ?: 0;
    0  1  ?  1  1: 0;
    0  0  0  0  ?: 0;
    0  0  ?  1  0: 0;
  endtable
endprimitive

primitive ADHCM2R_udp_0(CO,A, NCI);
  output CO;
  input A, NCI;
  table
  //A, NCI: CO
    1  0: 1;
    0  ?: 0;
    ?  1: 0;
  endtable
endprimitive

primitive ADHCM2R_udp_1(S,A, NCI);
  output S;
  input A, NCI;
  table
  //A, NCI: S
    1  1: 1;
    0  0: 1;
    1  0: 0;
    0  1: 0;
  endtable
endprimitive

primitive ADHCSCM2R_udp_0(S,A, CS, NCI);
  output S;
  input A, CS, NCI;
  table
  //A, CS, NCI: S
    1  0  ?: 1;
    1  ?  1: 1;
    0  1  0: 1;
    1  1  0: 0;
    0  0  ?: 0;
    0  ?  1: 0;
  endtable
endprimitive

primitive ADHCSOM2R_udp_0(S,A, CI, CS);
  output S;
  input A, CI, CS;
  table
  //A, CI, CS: S
    1  0  ?: 1;
    1  ?  0: 1;
    0  1  1: 1;
    1  1  1: 0;
    0  0  ?: 0;
    0  ?  0: 0;
  endtable
endprimitive

primitive ADHM1RA_udp_0(CO,A, B);
  output CO;
  input A, B;
  table
  //A, B: CO
    1  1: 1;
    0  ?: 0;
    ?  0: 0;
  endtable
endprimitive

primitive ADHM1RA_udp_1(S,A, B);
  output S;
  input A, B;
  table
  //A, B: S
    1  0: 1;
    0  1: 1;
    1  1: 0;
    0  0: 0;
  endtable
endprimitive

primitive AN3M0R_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    1  1  1: 1;
    0  ?  ?: 0;
    ?  0  ?: 0;
    ?  ?  0: 0;
  endtable
endprimitive

primitive AN4M0R_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  1  1  1: 1;
    0  ?  ?  ?: 0;
    ?  0  ?  ?: 0;
    ?  ?  0  ?: 0;
    ?  ?  ?  0: 0;
  endtable
endprimitive

primitive AO211M1RA_udp_0(Z,A1, A2, B, C);
  output Z;
  input A1, A2, B, C;
  table
  //A1, A2, B, C: Z
    1  1  ?  ?: 1;
    ?  ?  1  ?: 1;
    ?  ?  ?  1: 1;
    0  ?  0  0: 0;
    ?  0  0  0: 0;
  endtable
endprimitive

primitive AO21M0RA_udp_0(Z,A1, A2, B);
  output Z;
  input A1, A2, B;
  table
  //A1, A2, B: Z
    1  1  ?: 1;
    ?  ?  1: 1;
    0  ?  0: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive AO221M1RA_udp_0(Z,A1, A2, B1, B2, C);
  output Z;
  input A1, A2, B1, B2, C;
  table
  //A1, A2, B1, B2, C: Z
    1  1  ?  ?  ?: 1;
    ?  ?  1  1  ?: 1;
    ?  ?  ?  ?  1: 1;
    0  ?  0  ?  0: 0;
    0  ?  ?  0  0: 0;
    ?  0  0  ?  0: 0;
    ?  0  ?  0  0: 0;
  endtable
endprimitive

primitive AO222M1RA_udp_0(Z,A1, A2, B1, B2, C1, C2);
  output Z;
  input A1, A2, B1, B2, C1, C2;
  table
  //A1, A2, B1, B2, C1, C2: Z
    1  1  ?  ?  ?  ?: 1;
    ?  ?  1  1  ?  ?: 1;
    ?  ?  ?  ?  1  1: 1;
    0  ?  0  ?  0  ?: 0;
    0  ?  0  ?  ?  0: 0;
    0  ?  ?  0  0  ?: 0;
    0  ?  ?  0  ?  0: 0;
    ?  0  0  ?  0  ?: 0;
    ?  0  0  ?  ?  0: 0;
    ?  0  ?  0  0  ?: 0;
    ?  0  ?  0  ?  0: 0;
  endtable
endprimitive

primitive AO22B10M0R_udp_0(Z,A1, NA2, B1, B2);
  output Z;
  input A1, NA2, B1, B2;
  table
  //A1, NA2, B1, B2: Z
    1  0  ?  ?: 1;
    ?  ?  1  1: 1;
    0  ?  0  ?: 0;
    0  ?  ?  0: 0;
    ?  1  0  ?: 0;
    ?  1  ?  0: 0;
  endtable
endprimitive

primitive AO22B11M0R_udp_0(Z,A1, NA2, B1, NB2);
  output Z;
  input A1, NA2, B1, NB2;
  table
  //A1, NA2, B1, NB2: Z
    1  0  ?  ?: 1;
    ?  ?  1  0: 1;
    0  ?  0  ?: 0;
    0  ?  ?  1: 0;
    ?  1  0  ?: 0;
    ?  1  ?  1: 0;
  endtable
endprimitive

primitive AO22M0RA_udp_0(Z,A1, A2, B1, B2);
  output Z;
  input A1, A2, B1, B2;
  table
  //A1, A2, B1, B2: Z
    1  1  ?  ?: 1;
    ?  ?  1  1: 1;
    0  ?  0  ?: 0;
    0  ?  ?  0: 0;
    ?  0  0  ?: 0;
    ?  0  ?  0: 0;
  endtable
endprimitive

primitive AO31M1RA_udp_0(Z,A1, A2, A3, B);
  output Z;
  input A1, A2, A3, B;
  table
  //A1, A2, A3, B: Z
    1  1  1  ?: 1;
    ?  ?  ?  1: 1;
    0  ?  ?  0: 0;
    ?  0  ?  0: 0;
    ?  ?  0  0: 0;
  endtable
endprimitive

primitive AO32M1RA_udp_0(Z,A1, A2, A3, B1, B2);
  output Z;
  input A1, A2, A3, B1, B2;
  table
  //A1, A2, A3, B1, B2: Z
    1  1  1  ?  ?: 1;
    ?  ?  ?  1  1: 1;
    0  ?  ?  0  ?: 0;
    0  ?  ?  ?  0: 0;
    ?  0  ?  0  ?: 0;
    ?  0  ?  ?  0: 0;
    ?  ?  0  0  ?: 0;
    ?  ?  0  ?  0: 0;
  endtable
endprimitive

primitive AO33M1RA_udp_0(Z,A1, A2, A3, B1, B2, B3);
  output Z;
  input A1, A2, A3, B1, B2, B3;
  table
  //A1, A2, A3, B1, B2, B3: Z
    1  1  1  ?  ?  ?: 1;
    ?  ?  ?  1  1  1: 1;
    0  ?  ?  0  ?  ?: 0;
    0  ?  ?  ?  0  ?: 0;
    0  ?  ?  ?  ?  0: 0;
    ?  0  ?  0  ?  ?: 0;
    ?  0  ?  ?  0  ?: 0;
    ?  0  ?  ?  ?  0: 0;
    ?  ?  0  0  ?  ?: 0;
    ?  ?  0  ?  0  ?: 0;
    ?  ?  0  ?  ?  0: 0;
  endtable
endprimitive

primitive AOI211M0R_udp_0(Z,A1, B, C, A2);
  output Z;
  input A1, B, C, A2;
  table
  //A1, B, C, A2: Z
    0  0  0  ?: 1;
    ?  0  0  0: 1;
    1  ?  ?  1: 0;
    ?  1  ?  ?: 0;
    ?  ?  1  ?: 0;
  endtable
endprimitive

primitive AOI21B01M0R_udp_0(Z,A1, NB, A2);
  output Z;
  input A1, NB, A2;
  table
  //A1, NB, A2: Z
    0  1  ?: 1;
    ?  1  0: 1;
    1  ?  1: 0;
    ?  0  ?: 0;
  endtable
endprimitive

primitive AOI21B10M0R_udp_0(Z,A1, B, NA2);
  output Z;
  input A1, B, NA2;
  table
  //A1, B, NA2: Z
    0  0  ?: 1;
    ?  0  1: 1;
    1  ?  0: 0;
    ?  1  ?: 0;
  endtable
endprimitive

primitive AOI21B20M0R_udp_0(Z,B, NA1, NA2);
  output Z;
  input B, NA1, NA2;
  table
  //B, NA1, NA2: Z
    0  1  ?: 1;
    0  ?  1: 1;
    1  ?  ?: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive AOI21M0R_udp_0(Z,A1, B, A2);
  output Z;
  input A1, B, A2;
  table
  //A1, B, A2: Z
    0  0  ?: 1;
    ?  0  0: 1;
    1  ?  1: 0;
    ?  1  ?: 0;
  endtable
endprimitive

primitive AOI221M0R_udp_0(Z,A1, B1, C, B2, A2);
  output Z;
  input A1, B1, C, B2, A2;
  table
  //A1, B1, C, B2, A2: Z
    0  0  0  ?  ?: 1;
    0  ?  0  0  ?: 1;
    ?  0  0  ?  0: 1;
    ?  ?  0  0  0: 1;
    1  ?  ?  ?  1: 0;
    ?  1  ?  1  ?: 0;
    ?  ?  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI222M0RA_udp_0(Z,A1, B1, C1, C2, B2, A2);
  output Z;
  input A1, B1, C1, C2, B2, A2;
  table
  //A1, B1, C1, C2, B2, A2: Z
    0  0  0  ?  ?  ?: 1;
    0  0  ?  0  ?  ?: 1;
    0  ?  0  ?  0  ?: 1;
    0  ?  ?  0  0  ?: 1;
    ?  0  0  ?  ?  0: 1;
    ?  0  ?  0  ?  0: 1;
    ?  ?  0  ?  0  0: 1;
    ?  ?  ?  0  0  0: 1;
    1  ?  ?  ?  ?  1: 0;
    ?  1  ?  ?  1  ?: 0;
    ?  ?  1  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI22B20M0R_udp_0(Z,B1, NA1, NA2, B2);
  output Z;
  input B1, NA1, NA2, B2;
  table
  //B1, NA1, NA2, B2: Z
    0  1  ?  ?: 1;
    0  ?  1  ?: 1;
    ?  1  ?  0: 1;
    ?  ?  1  0: 1;
    1  ?  ?  1: 0;
    ?  0  0  ?: 0;
  endtable
endprimitive

primitive AOI22M0R_udp_0(Z,A1, B1, B2, A2);
  output Z;
  input A1, B1, B2, A2;
  table
  //A1, B1, B2, A2: Z
    0  0  ?  ?: 1;
    0  ?  0  ?: 1;
    ?  0  ?  0: 1;
    ?  ?  0  0: 1;
    1  ?  ?  1: 0;
    ?  1  1  ?: 0;
  endtable
endprimitive

primitive AOI31M0R_udp_0(Z,A1, B, A2, A3);
  output Z;
  input A1, B, A2, A3;
  table
  //A1, B, A2, A3: Z
    0  0  ?  ?: 1;
    ?  0  0  ?: 1;
    ?  0  ?  0: 1;
    1  ?  1  1: 0;
    ?  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI32M0R_udp_0(Z,A1, B1, B2, A2, A3);
  output Z;
  input A1, B1, B2, A2, A3;
  table
  //A1, B1, B2, A2, A3: Z
    0  0  ?  ?  ?: 1;
    0  ?  0  ?  ?: 1;
    ?  0  ?  0  ?: 1;
    ?  ?  0  0  ?: 1;
    ?  0  ?  ?  0: 1;
    ?  ?  0  ?  0: 1;
    1  ?  ?  1  1: 0;
    ?  1  1  ?  ?: 0;
  endtable
endprimitive

primitive AOI33M0R_udp_0(Z,A1, B1, B2, B3, A2, A3);
  output Z;
  input A1, B1, B2, B3, A2, A3;
  table
  //A1, B1, B2, B3, A2, A3: Z
    0  0  ?  ?  ?  ?: 1;
    0  ?  0  ?  ?  ?: 1;
    0  ?  ?  0  ?  ?: 1;
    ?  0  ?  ?  0  ?: 1;
    ?  ?  0  ?  0  ?: 1;
    ?  ?  ?  0  0  ?: 1;
    ?  0  ?  ?  ?  0: 1;
    ?  ?  0  ?  ?  0: 1;
    ?  ?  ?  0  ?  0: 1;
    1  ?  ?  ?  1  1: 0;
    ?  1  1  1  ?  ?: 0;
  endtable
endprimitive

primitive BEM2RA_udp_0(OA1,M0, M1, M2);
  output OA1;
  input M0, M1, M2;
  table
  //M0, M1, M2: OA1
    1  1  ?: 1;
    ?  ?  0: 1;
    0  ?  1: 0;
    ?  0  1: 0;
  endtable
endprimitive

primitive BEM2RA_udp_1(OA2,M0, M1, M2);
  output OA2;
  input M0, M1, M2;
  table
  //M0, M1, M2: OA2
    0  0  ?: 1;
    ?  ?  1: 1;
    1  ?  0: 0;
    ?  1  0: 0;
  endtable
endprimitive

primitive BEMXBM2R_udp_0(PB,M0, OA1, Z, OA2, M1);
  output PB;
  input M0, OA1, Z, OA2, M1;
  table
  //M0, OA1, Z, OA2, M1: PB
    1  1  1  ?  ?: 1;
    0  ?  1  1  ?: 1;
    ?  1  0  ?  1: 1;
    ?  ?  0  1  0: 1;
    ?  1  ?  1  ?: 1;
    1  0  1  ?  ?: 0;
    0  ?  1  0  ?: 0;
    ?  0  0  ?  1: 0;
    ?  ?  0  0  0: 0;
    ?  0  ?  0  ?: 0;
  endtable
endprimitive

primitive BEMXM2RA_udp_0(P,M0, OA1, Z, OA2, M1);
  output P;
  input M0, OA1, Z, OA2, M1;
  table
  //M0, OA1, Z, OA2, M1: P
    1  0  1  ?  ?: 1;
    0  ?  1  0  ?: 1;
    ?  0  0  ?  1: 1;
    ?  ?  0  0  0: 1;
    ?  0  ?  0  ?: 1;
    1  1  1  ?  ?: 0;
    0  ?  1  1  ?: 0;
    ?  1  0  ?  1: 0;
    ?  ?  0  1  0: 0;
    ?  1  ?  1  ?: 0;
  endtable
endprimitive

primitive BUFTM0R_udp_0(MGM_WB_0,A, E);
  output MGM_WB_0;
  input A, E;
  table
  //A, E: MGM_WB_0
    1  1: 1;
    0  1: 0;
    ?  0: 1;   
  endtable
endprimitive

primitive CKMUX2M12R_udp_0(Z,A, S, B);
  output Z;
  input A, S, B;
  table
  //A, S, B: Z
    1  0  ?: 1;
    ?  1  1: 1;
    0  0  ?: 0;
    ?  1  0: 0;
    1  ?  1: 1;
    0  ?  0: 0;
  endtable
endprimitive

primitive DFEM1RA_udp_0(MGM_D,D, E, IQ);
  output MGM_D;
  input D, E, IQ;
  table
  //D, E, IQ: MGM_D
    1  1  ?: 1;
    1  ?  1: 1;
    ?  0  1: 1;
    0  1  ?: 0;
    0  ?  0: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive DFEQZRM1RA_udp_0(MGM_D,D, E, RB, IQ);
  output MGM_D;
  input D, E, RB, IQ;
  table
  //D, E, RB, IQ: MGM_D
    1  1  1  ?: 1;
    1  ?  1  1: 1;
    ?  0  1  1: 1;
    0  1  ?  ?: 0;
    0  ?  ?  0: 0;
    ?  0  ?  0: 0;
    ?  ?  0  ?: 0;
  endtable
endprimitive

primitive DFMM1RA_udp_0(MGM_D,D1, S, D2);
  output MGM_D;
  input D1, S, D2;
  table
  //D1, S, D2: MGM_D
    1  1  ?: 1;
    ?  0  1: 1;
    0  1  ?: 0;
    ?  0  0: 0;
    1  ?  1: 1;
    0  ?  0: 0;
  endtable
endprimitive

primitive DFQZRSM1RA_udp_0(MGM_D,D, RB, SB);
  output MGM_D;
  input D, RB, SB;
  table
  //D, RB, SB: MGM_D
    1  1  ?: 1;
    ?  1  0: 1;
    0  ?  1: 0;
    ?  0  ?: 0;
  endtable
endprimitive

primitive DFQZSM1RA_udp_0(MGM_D,D, SB);
  output MGM_D;
  input D, SB;
  table
  //D, SB: MGM_D
    1  ?: 1;
    ?  0: 1;
    0  1: 0;
  endtable
endprimitive

primitive LAGCECSM12RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;


endtable
endprimitive

primitive LAGCECSM16RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;


endtable
endprimitive

primitive LAGCECSM24RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM2RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM32RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM40RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM48RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM4RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM6RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCECSM8RA_statetable_ENL(ENL,CKB,E,SE);
output ENL ;
reg ENL;
input CKB,E,SE; 
table 
//CKB E SE : ENL : ENL
  1  0  0   : ?   : 0;
  1  ?  1   : ?   : 1;
  1  1  ?   : ?   : 1;
  0  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM12R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM16R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM20R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM2R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM3R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM4R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM6R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEM8R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM12R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM12R_udp_0(GCK,CK, ENL, SE);
  output GCK;
  input CK, ENL, SE;
  table
  //CK, ENL, SE: GCK
    1  1  ?: 1;
    1  ?  1: 1;
    0  ?  ?: 0;
    ?  0  0: 0;
  endtable
endprimitive

primitive LAGCEPM16R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM20R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM2R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM3R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM4R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM6R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPM8R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM12R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM16R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM20R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM2R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM3R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM4R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM6R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCEPOM8R_statetable_ENL(ENL,CK,E);
output ENL ;
reg ENL;
input CK,E; 
table 
//CK E : ENL : ENL
  0  0   : ?   : 0;
  0  1   : ?   : 1;
  1  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM12RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM16RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM24RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM2RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM32RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM40RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM48RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM4RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM6RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESM8RA_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM12R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM16R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM20R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM2R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM3R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM4R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM6R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive LAGCESOM8R_statetable_ENL(ENL,CK,E,SE);
output ENL ;
reg ENL;
input CK,E,SE; 
table 
//CK E SE : ENL : ENL
  0  0  0   : ?   : 0;
  0  ?  1   : ?   : 1;
  0  1  ?   : ?   : 1;
  1  ?  ?   : ?   : -;

endtable
endprimitive

primitive MAOI2223M1RA_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    0  0  0  ?: 1;
    0  ?  ?  0: 1;
    ?  0  ?  0: 1;
    ?  ?  0  0: 1;
    1  1  1  ?: 0;
    1  ?  ?  1: 0;
    ?  1  ?  1: 0;
    ?  ?  1  1: 0;
  endtable
endprimitive

primitive MGM_H_IQ_LATCH_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  Q  :  Q 
  ?  ?  0  *  ?  :  ?  :  -;  // No change CK=0
  ?  0  1  0  ?  :  ?  :  0;  // Latch 0 
  ?  0  *  0  ?  :  0  :  0;  // reduce pessimism when D=0
  1  0  ?  ?  ?  :  ?  :  0;  // clear
  0  ?  1  1  ?  :  ?  :  1;  // Latch 1
  0  ?  *  1  ?  :  1  :  1;  // reduce pessimism when D=1
  ?  1  ?  ?  ?  :  ?  :  1;  // Preset P dominate C
  *  0  0  ?  ?  :  0  :  0;   // reduce clear pessimism
  *  0  ?  0  ?  :  0  :  0;   // reduce clear pessimism
  0  *  0  ?  ?  :  1  :  1;   // reduce preset pessimism
  0  *  ?  1  ?  :  1  :  1;   // reduce preset pessimism

//  ?  ?  ?  ?  *  :  ?  :  x;  // notifier
                  
endtable
endprimitive

primitive MGM_H_IQN_FF_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  QN  :  QN 
  ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  1;  // CK in 0
  ?  0  p  0  ?  :  1  :  1;  // reduce pessimism D=0
  1  ?  ?  ?  ?  :  ?  :  1;  // clear: C dominate P
  0  ?  r  1  ?  :  ?  :  0;  // CK in 1
  0  ?  p  1  ?  :  0  :  0;  // reduce pessimism D=1
  0  1  ?  ?  ?  :  ?  :  0;  // preset
  ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
  *  0  b  ?  ?  :  1  :  1;  // reduce clear pessimism
  *  0  x  0  ?  :  1  :  1;  // reduce clear pessimism
  0  *  b  ?  ?  :  0  :  0;  // reduce preset pessimism
  0  *  x  1  ?  :  0  :  0;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_IQ_FF_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//  C  P  CK  D  N :  Q  :  Q 
    ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
    ?  0  r  0  ?  :  ?  :  0;  // CK in 0
    ?  0  p  0  ?  :  0  :  0;  // reduce pessimism D=0
    1  ?  ?  ?  ?  :  ?  :  0;  // clear: C dominate P
    0  ?  r  1  ?  :  ?  :  1;  // CK in 1
    0  ?  p  1  ?  :  1  :  1;  // reduce pessimism D=1
    0  1  ?  ?  ?  :  ?  :  1;  // preset
    ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
    *  0  b  ?  ?  :  0  :  0;  // reduce clear pessimism
    *  0  x  0  ?  :  0  :  0;  // reduce clear pessimism
    0  *  b  ?  ?  :  1  :  1;  // reduce preset pessimism
    0  *  x  1  ?  :  1  :  1;  // reduce preset pessimism
//  ?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_IQ_LATCH_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//  C  P  CK  D  N :  Q  :  Q 
    ?  ?  0  *  ?  :  ?  :  -;   // No change CK=0
    ?  0  1  0  ?  :  ?  :  0;   // Latch 0
    ?  0  *  0  ?  :  0  :  0;   // reduce pessimism when D=0
    1  ?  ?  ?  ?  :  ?  :  0;   // Clear : C dominate P
    0  ?  1  1  ?  :  ?  :  1;   // Latch 1
    0  ?  *  1  ?  :  1  :  1;   // reduce pessimism when D=1
    0  1  ?  ?  ?  :  ?  :  1;   // Preset
    *  0  0  ?  ?  :  0  :  0;   // reduce clear pessimism
    *  0  ?  0  ?  :  0  :  0;   // reduce clear pessimism
    0  *  0  ?  ?  :  1  :  1;   // reduce preset pessimism
    0  *  ?  1  ?  :  1  :  1;   // reduce preset pessimism
//  ?  ?  ?  ?  *  :  ?  :  x;   // notifier
                  
endtable
endprimitive

primitive MGM_IQN_FF_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  QN  :  QN 
  ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  1;  // CK in 0
  ?  0  p  0  ?  :  1  :  1;  // reduce pessimism D=0
  1  ?  ?  ?  ?  :  ?  :  1;  // clear: C dominate P
  0  ?  r  1  ?  :  ?  :  0;  // CK in 1
  0  ?  p  1  ?  :  0  :  0;  // reduce pessimism D=1
  0  1  ?  ?  ?  :  ?  :  0;  // preset
  ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
  *  0  b  ?  ?  :  1  :  1;  // reduce clear pessimism
  *  0  x  0  ?  :  1  :  1;  // reduce clear pessimism
  0  *  b  ?  ?  :  0  :  0;  // reduce preset pessimism
  0  *  x  1  ?  :  0  :  0;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_IQN_LATCH_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N : QN : QN 
  ?  ?  0  *  ?  :  ?  :  -;  // No change CK=0
  ?  0  1  0  ?  :  ?  :  1;  // Latch 0
  ?  0  *  0  ?  :  1  :  1;  // reduce pessimism when D=0
  1  ?  ?  ?  ?  :  ?  :  1;  // Clear : C dominate P
  0  ?  1  1  ?  :  ?  :  0;  // Latch 1
  0  ?  *  1  ?  :  0  :  0;  // reduce pessimism when D=1
  0  1  ?  ?  ?  :  ?  :  0;  // Preset
  *  0  0  ?  ?  :  1  :  1;   // reduce clear pessimism
  *  0  ?  0  ?  :  1  :  1;   // reduce clear pessimism
  0  *  0  ?  ?  :  0  :  0;   // reduce preset pessimism
  0  *  ?  1  ?  :  0  :  0;   // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;   // notifier
                  
endtable
endprimitive

primitive MGM_L_IQ_FF_UDP(Q,C,P,CK,D,N);
output Q;
reg Q;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  Q  :  Q 
  ?  ?  n  ?  ?  :  ?  :  -;  // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  0;  // CK in 0
  ?  0  p  0  ?  :  0  :  0;  // reduce pessimism D=0
  1  ?  ?  ?  ?  :  ?  :  0;  // clear: C dominate P
  0  ?  r  1  ?  :  ?  :  1;  // CK in 1
  0  ?  p  1  ?  :  1  :  1;  // reduce pessimism D=1
  0  1  ?  ?  ?  :  ?  :  1;  // preset
  ?  ?  b  *  ?  :  ?  :  -;  // ignore D change on steady CK
  *  0  b  ?  ?  :  0  :  0;  // reduce clear pessimism
  *  0  x  0  ?  :  0  :  0;  // reduce clear pessimism
  0  *  b  ?  ?  :  1  :  1;  // reduce preset pessimism
  0  *  x  1  ?  :  1  :  1;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x;  // notifier change
                  
endtable
endprimitive

primitive MGM_L_IQN_FF_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N :  QN  :  QN 
  ?  ?  n  ?  ?  :  ?  :  -; // no changes on neg CK
  ?  0  r  0  ?  :  ?  :  1; // CK in 0
  ?  0  p  0  ?  :  1  :  1; // reduce pessimism D=0
  1  0  ?  ?  ?  :  ?  :  1; // clear
  0  ?  r  1  ?  :  ?  :  0; // CK in 1
  0  ?  p  1  ?  :  0  :  0; // reduce pessimism D=1
  ?  1  ?  ?  ?  :  ?  :  0; // preset P dominate C
  ?  ?  b  *  ?  :  ?  :  -; // ignore D change on steady CK : add
  *  0  b  ?  ?  :  1  :  1;  // reduce clear pessimism
  *  0  x  0  ?  :  1  :  1;  // reduce clear pessimism
  0  *  b  ?  ?  :  0  :  0;  // reduce preset pessimism
  0  *  x  1  ?  :  0  :  0;  // reduce preset pessimism
//?  ?  ?  ?  *  :  ?  :  x; // notifier change
                  
endtable
endprimitive

primitive MGM_L_IQN_LATCH_UDP(QN,C,P,CK,D,N);
output QN;
reg QN;
input C,P,CK,D,N; 
table 
//C  P  CK  D  N : QN : QN 
  ?  ?  0  *  ?  :  ?  :  -;  // No change CK=0
  ?  0  1  0  ?  :  ?  :  1;  // Latch 0
  ?  0  *  0  ?  :  1  :  1;  // reduce pessimism when D=0
  1  0  ?  ?  ?  :  ?  :  1;  // clear
  0  ?  1  1  ?  :  ?  :  0;  // Latch 1
  0  ?  *  1  ?  :  0  :  0;  // reduce pessimism when D=1
  ?  1  ?  ?  ?  :  ?  :  0;  // Preset P dominate C
  *  0  0  ?  ?  :  1  :  1;   // reduce clear pessimism
  *  0  ?  0  ?  :  1  :  1;   // reduce clear pessimism
  0  *  0  ?  ?  :  0  :  0;   // reduce preset pessimism
  0  *  ?  1  ?  :  0  :  0;   // reduce preset pessimism

//  ?  ?  ?  ?  *  :  ?  :  x;  // notifier
                  
endtable
endprimitive

primitive MOAI22M1RA_udp_0(Z,A1, A2, B1, B2);
  output Z;
  input A1, A2, B1, B2;
  table
  //A1, A2, B1, B2: Z
    0  0  ?  ?: 1;
    ?  ?  1  1: 1;
    1  ?  0  ?: 0;
    1  ?  ?  0: 0;
    ?  1  0  ?: 0;
    ?  1  ?  0: 0;
  endtable
endprimitive

primitive MUX3M0RA_udp_0(Z,A, S0, S1, B, C);
  output Z;
  input A, S0, S1, B, C;
  table
  //A, S0, S1, B, C: Z
    1  0  0  ?  ?: 1;
    ?  1  0  1  ?: 1;
    ?  ?  1  ?  1: 1;
    0  0  0  ?  ?: 0;
    ?  1  0  0  ?: 0;
    ?  ?  1  ?  0: 0;
    1  ?  0  1  ?: 1;
    ?  1  ?  1  1: 1;
    1  0  ?  ?  1: 1;
    1  ?  ?  1  1: 1;
    0  ?  0  0  ?: 0;
    ?  1  ?  0  0: 0;
    0  0  ?  ?  0: 0;
    0  ?  ?  0  0: 0;
  endtable
endprimitive

primitive MUX4M0RA_udp_0(Z,A, S0, S1, B, C, D);
  output Z;
  input A, S0, S1, B, C, D;
  table
  //A, S0, S1, B, C, D: Z
    1  0  0  ?  ?  ?: 1;
    ?  1  0  1  ?  ?: 1;
    ?  0  1  ?  1  ?: 1;
    ?  1  1  ?  ?  1: 1;
    0  0  0  ?  ?  ?: 0;
    ?  1  0  0  ?  ?: 0;
    ?  0  1  ?  0  ?: 0;
    ?  1  1  ?  ?  0: 0;
    1  ?  0  1  ?  ?: 1;
    ?  ?  1  ?  1  1: 1;
    1  0  ?  ?  1  ?: 1;
    ?  1  ?  1  ?  1: 1;
    1  ?  ?  1  1  1: 1;
    0  ?  0  0  ?  ?: 0;
    ?  ?  1  ?  0  0: 0;
    0  0  ?  ?  0  ?: 0;
    ?  1  ?  0  ?  0: 0;
    0  ?  ?  0  0  0: 0;
  endtable
endprimitive

primitive MXB2M0RA_udp_0(Z,A, S, B);
  output Z;
  input A, S, B;
  table
  //A, S, B: Z
    0  0  ?: 1;
    ?  1  0: 1;
    1  0  ?: 0;
    ?  1  1: 0;
    1  ?  1: 0;
    0  ?  0: 1;
  endtable
endprimitive

primitive MXB3M0RA_udp_0(Z,A, S0, S1, B, C);
  output Z;
  input A, S0, S1, B, C;
  table
  //A, S0, S1, B, C: Z
    0  0  0  ?  ?: 1;
    ?  1  0  0  ?: 1;
    ?  ?  1  ?  0: 1;
    1  0  0  ?  ?: 0;
    ?  1  0  1  ?: 0;
    ?  ?  1  ?  1: 0;
    1  ?  0  1  ?: 0;
    ?  1  ?  1  1: 0;
    1  0  ?  ?  1: 0;
    1  ?  ?  1  1: 0;
    0  ?  0  0  ?: 1;
    ?  1  ?  0  0: 1;
    0  0  ?  ?  0: 1;
    0  ?  ?  0  0: 1;
  endtable
endprimitive

primitive MXB4M0RA_udp_0(Z,A, S0, S1, B, C, D);
  output Z;
  input A, S0, S1, B, C, D;
  table
  //A, S0, S1, B, C, D: Z
    0  0  0  ?  ?  ?: 1;
    ?  1  0  0  ?  ?: 1;
    ?  0  1  ?  0  ?: 1;
    ?  1  1  ?  ?  0: 1;
    1  0  0  ?  ?  ?: 0;
    ?  1  0  1  ?  ?: 0;
    ?  0  1  ?  1  ?: 0;
    ?  1  1  ?  ?  1: 0;
    1  ?  0  1  ?  ?: 0;
    ?  ?  1  ?  1  1: 0;
    1  0  ?  ?  1  ?: 0;
    ?  1  ?  1  ?  1: 0;
    1  ?  ?  1  1  1: 0;
    0  ?  0  0  ?  ?: 1;
    ?  ?  1  ?  0  0: 1;
    0  0  ?  ?  0  ?: 1;
    ?  1  ?  0  ?  0: 1;
    0  ?  ?  0  0  0: 1;
  endtable
endprimitive

primitive ND2B1M0R_udp_0(Z,B, NA);
  output Z;
  input B, NA;
  table
  //B, NA: Z
    0  ?: 1;
    ?  1: 1;
    1  0: 0;
  endtable
endprimitive

primitive ND3B1M0R_udp_0(Z,B, C, NA);
  output Z;
  input B, C, NA;
  table
  //B, C, NA: Z
    0  ?  ?: 1;
    ?  0  ?: 1;
    ?  ?  1: 1;
    1  1  0: 0;
  endtable
endprimitive

primitive ND3M0R_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    0  ?  ?: 1;
    ?  0  ?: 1;
    ?  ?  0: 1;
    1  1  1: 0;
  endtable
endprimitive

primitive ND4B1M0R_udp_0(Z,B, C, D, NA);
  output Z;
  input B, C, D, NA;
  table
  //B, C, D, NA: Z
    0  ?  ?  ?: 1;
    ?  0  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  1: 1;
    1  1  1  0: 0;
  endtable
endprimitive

primitive ND4B2M0R_udp_0(Z,C, D, NA, NB);
  output Z;
  input C, D, NA, NB;
  table
  //C, D, NA, NB: Z
    0  ?  ?  ?: 1;
    ?  0  ?  ?: 1;
    ?  ?  1  ?: 1;
    ?  ?  ?  1: 1;
    1  1  0  0: 0;
  endtable
endprimitive

primitive ND4M0R_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    0  ?  ?  ?: 1;
    ?  0  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  0: 1;
    1  1  1  1: 0;
  endtable
endprimitive

primitive NR2B1M0R_udp_0(Z,B, NA);
  output Z;
  input B, NA;
  table
  //B, NA: Z
    0  1: 1;
    1  ?: 0;
    ?  0: 0;
  endtable
endprimitive

primitive NR3B1M0R_udp_0(Z,B, C, NA);
  output Z;
  input B, C, NA;
  table
  //B, C, NA: Z
    0  0  1: 1;
    1  ?  ?: 0;
    ?  1  ?: 0;
    ?  ?  0: 0;
  endtable
endprimitive

primitive NR3M0R_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    0  0  0: 1;
    1  ?  ?: 0;
    ?  1  ?: 0;
    ?  ?  1: 0;
  endtable
endprimitive

primitive NR4B1M0R_udp_0(Z,B, C, D, NA);
  output Z;
  input B, C, D, NA;
  table
  //B, C, D, NA: Z
    0  0  0  1: 1;
    1  ?  ?  ?: 0;
    ?  1  ?  ?: 0;
    ?  ?  1  ?: 0;
    ?  ?  ?  0: 0;
  endtable
endprimitive

primitive NR4B2M0R_udp_0(Z,C, D, NA, NB);
  output Z;
  input C, D, NA, NB;
  table
  //C, D, NA, NB: Z
    0  0  1  1: 1;
    1  ?  ?  ?: 0;
    ?  1  ?  ?: 0;
    ?  ?  0  ?: 0;
    ?  ?  ?  0: 0;
  endtable
endprimitive

primitive NR4M0R_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    0  0  0  0: 1;
    1  ?  ?  ?: 0;
    ?  1  ?  ?: 0;
    ?  ?  1  ?: 0;
    ?  ?  ?  1: 0;
  endtable
endprimitive

primitive OA211M12RA_udp_0(Z,A1, B, C, A2);
  output Z;
  input A1, B, C, A2;
  table
  //A1, B, C, A2: Z
    1  1  1  ?: 1;
    ?  1  1  1: 1;
    0  ?  ?  0: 0;
    ?  0  ?  ?: 0;
    ?  ?  0  ?: 0;
  endtable
endprimitive

primitive OA21M0RA_udp_0(Z,A1, B, A2);
  output Z;
  input A1, B, A2;
  table
  //A1, B, A2: Z
    1  1  ?: 1;
    ?  1  1: 1;
    0  ?  0: 0;
    ?  0  ?: 0;
  endtable
endprimitive

primitive OA221M1RA_udp_0(Z,A1, B1, C, B2, A2);
  output Z;
  input A1, B1, C, B2, A2;
  table
  //A1, B1, C, B2, A2: Z
    1  1  1  ?  ?: 1;
    1  ?  1  1  ?: 1;
    ?  1  1  ?  1: 1;
    ?  ?  1  1  1: 1;
    0  ?  ?  ?  0: 0;
    ?  0  ?  0  ?: 0;
    ?  ?  0  ?  ?: 0;
  endtable
endprimitive

primitive OA222M1RA_udp_0(Z,A1, B1, C1, C2, B2, A2);
  output Z;
  input A1, B1, C1, C2, B2, A2;
  table
  //A1, B1, C1, C2, B2, A2: Z
    1  1  1  ?  ?  ?: 1;
    1  1  ?  1  ?  ?: 1;
    1  ?  1  ?  1  ?: 1;
    1  ?  ?  1  1  ?: 1;
    ?  1  1  ?  ?  1: 1;
    ?  1  ?  1  ?  1: 1;
    ?  ?  1  ?  1  1: 1;
    ?  ?  ?  1  1  1: 1;
    0  ?  ?  ?  ?  0: 0;
    ?  0  ?  ?  0  ?: 0;
    ?  ?  0  0  ?  ?: 0;
  endtable
endprimitive

primitive OA22M0R_udp_0(Z,A1, B1, B2, A2);
  output Z;
  input A1, B1, B2, A2;
  table
  //A1, B1, B2, A2: Z
    1  1  ?  ?: 1;
    1  ?  1  ?: 1;
    ?  1  ?  1: 1;
    ?  ?  1  1: 1;
    0  ?  ?  0: 0;
    ?  0  0  ?: 0;
  endtable
endprimitive

primitive OA31M1RA_udp_0(Z,A1, B, A2, A3);
  output Z;
  input A1, B, A2, A3;
  table
  //A1, B, A2, A3: Z
    1  1  ?  ?: 1;
    ?  1  1  ?: 1;
    ?  1  ?  1: 1;
    0  ?  0  0: 0;
    ?  0  ?  ?: 0;
  endtable
endprimitive

primitive OA32M1RA_udp_0(Z,A1, B1, B2, A2, A3);
  output Z;
  input A1, B1, B2, A2, A3;
  table
  //A1, B1, B2, A2, A3: Z
    1  1  ?  ?  ?: 1;
    1  ?  1  ?  ?: 1;
    ?  1  ?  1  ?: 1;
    ?  ?  1  1  ?: 1;
    ?  1  ?  ?  1: 1;
    ?  ?  1  ?  1: 1;
    0  ?  ?  0  0: 0;
    ?  0  0  ?  ?: 0;
  endtable
endprimitive

primitive OA33M1RA_udp_0(Z,A1, B1, B2, B3, A2, A3);
  output Z;
  input A1, B1, B2, B3, A2, A3;
  table
  //A1, B1, B2, B3, A2, A3: Z
    1  1  ?  ?  ?  ?: 1;
    1  ?  1  ?  ?  ?: 1;
    1  ?  ?  1  ?  ?: 1;
    ?  1  ?  ?  1  ?: 1;
    ?  ?  1  ?  1  ?: 1;
    ?  ?  ?  1  1  ?: 1;
    ?  1  ?  ?  ?  1: 1;
    ?  ?  1  ?  ?  1: 1;
    ?  ?  ?  1  ?  1: 1;
    0  ?  ?  ?  0  0: 0;
    ?  0  0  0  ?  ?: 0;
  endtable
endprimitive

primitive OAI211B100M0R_udp_0(Z,A1, NA2, B, C);
  output Z;
  input A1, NA2, B, C;
  table
  //A1, NA2, B, C: Z
    0  1  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  0: 1;
    1  ?  1  1: 0;
    ?  0  1  1: 0;
  endtable
endprimitive

primitive OAI211M0R_udp_0(Z,A1, A2, B, C);
  output Z;
  input A1, A2, B, C;
  table
  //A1, A2, B, C: Z
    0  0  ?  ?: 1;
    ?  ?  0  ?: 1;
    ?  ?  ?  0: 1;
    1  ?  1  1: 0;
    ?  1  1  1: 0;
  endtable
endprimitive

primitive OAI21B10M0R_udp_0(Z,A1, NA2, B);
  output Z;
  input A1, NA2, B;
  table
  //A1, NA2, B: Z
    0  1  ?: 1;
    ?  ?  0: 1;
    1  ?  1: 0;
    ?  0  1: 0;
  endtable
endprimitive

primitive OAI21B20M0R_udp_0(Z,B, NA1, NA2);
  output Z;
  input B, NA1, NA2;
  table
  //B, NA1, NA2: Z
    0  ?  ?: 1;
    ?  1  1: 1;
    1  0  ?: 0;
    1  ?  0: 0;
  endtable
endprimitive

primitive OAI21M0R_udp_0(Z,A1, A2, B);
  output Z;
  input A1, A2, B;
  table
  //A1, A2, B: Z
    0  0  ?: 1;
    ?  ?  0: 1;
    1  ?  1: 0;
    ?  1  1: 0;
  endtable
endprimitive

primitive OAI221M0R_udp_0(Z,A1, A2, B1, B2, C);
  output Z;
  input A1, A2, B1, B2, C;
  table
  //A1, A2, B1, B2, C: Z
    0  0  ?  ?  ?: 1;
    ?  ?  0  0  ?: 1;
    ?  ?  ?  ?  0: 1;
    1  ?  1  ?  1: 0;
    1  ?  ?  1  1: 0;
    ?  1  1  ?  1: 0;
    ?  1  ?  1  1: 0;
  endtable
endprimitive

primitive OAI222M0RA_udp_0(Z,A1, A2, B1, B2, C1, C2);
  output Z;
  input A1, A2, B1, B2, C1, C2;
  table
  //A1, A2, B1, B2, C1, C2: Z
    0  0  ?  ?  ?  ?: 1;
    ?  ?  0  0  ?  ?: 1;
    ?  ?  ?  ?  0  0: 1;
    1  ?  1  ?  1  ?: 0;
    1  ?  1  ?  ?  1: 0;
    1  ?  ?  1  1  ?: 0;
    1  ?  ?  1  ?  1: 0;
    ?  1  1  ?  1  ?: 0;
    ?  1  1  ?  ?  1: 0;
    ?  1  ?  1  1  ?: 0;
    ?  1  ?  1  ?  1: 0;
  endtable
endprimitive

primitive OAI22B10M0R_udp_0(Z,A1, NA2, B1, B2);
  output Z;
  input A1, NA2, B1, B2;
  table
  //A1, NA2, B1, B2: Z
    0  1  ?  ?: 1;
    ?  ?  0  0: 1;
    1  ?  1  ?: 0;
    1  ?  ?  1: 0;
    ?  0  1  ?: 0;
    ?  0  ?  1: 0;
  endtable
endprimitive

primitive OAI22M0R_udp_0(Z,A1, A2, B1, B2);
  output Z;
  input A1, A2, B1, B2;
  table
  //A1, A2, B1, B2: Z
    0  0  ?  ?: 1;
    ?  ?  0  0: 1;
    1  ?  1  ?: 0;
    1  ?  ?  1: 0;
    ?  1  1  ?: 0;
    ?  1  ?  1: 0;
  endtable
endprimitive

primitive OAI31M0R_udp_0(Z,A1, A2, A3, B);
  output Z;
  input A1, A2, A3, B;
  table
  //A1, A2, A3, B: Z
    0  0  0  ?: 1;
    ?  ?  ?  0: 1;
    1  ?  ?  1: 0;
    ?  1  ?  1: 0;
    ?  ?  1  1: 0;
  endtable
endprimitive

primitive OAI32M0R_udp_0(Z,A1, A2, A3, B1, B2);
  output Z;
  input A1, A2, A3, B1, B2;
  table
  //A1, A2, A3, B1, B2: Z
    0  0  0  ?  ?: 1;
    ?  ?  ?  0  0: 1;
    1  ?  ?  1  ?: 0;
    1  ?  ?  ?  1: 0;
    ?  1  ?  1  ?: 0;
    ?  1  ?  ?  1: 0;
    ?  ?  1  1  ?: 0;
    ?  ?  1  ?  1: 0;
  endtable
endprimitive

primitive OAI33M0R_udp_0(Z,A1, A2, A3, B1, B2, B3);
  output Z;
  input A1, A2, A3, B1, B2, B3;
  table
  //A1, A2, A3, B1, B2, B3: Z
    0  0  0  ?  ?  ?: 1;
    ?  ?  ?  0  0  0: 1;
    1  ?  ?  1  ?  ?: 0;
    1  ?  ?  ?  1  ?: 0;
    1  ?  ?  ?  ?  1: 0;
    ?  1  ?  1  ?  ?: 0;
    ?  1  ?  ?  1  ?: 0;
    ?  1  ?  ?  ?  1: 0;
    ?  ?  1  1  ?  ?: 0;
    ?  ?  1  ?  1  ?: 0;
    ?  ?  1  ?  ?  1: 0;
  endtable
endprimitive

primitive OR2M0R_udp_0(Z,A, B);
  output Z;
  input A, B;
  table
  //A, B: Z
    1  ?: 1;
    ?  1: 1;
    0  0: 0;
  endtable
endprimitive

primitive OR3M0R_udp_0(Z,A, B, C);
  output Z;
  input A, B, C;
  table
  //A, B, C: Z
    1  ?  ?: 1;
    ?  1  ?: 1;
    ?  ?  1: 1;
    0  0  0: 0;
  endtable
endprimitive

primitive OR4M0R_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  ?  ?  ?: 1;
    ?  1  ?  ?: 1;
    ?  ?  1  ?: 1;
    ?  ?  ?  1: 1;
    0  0  0  0: 0;
  endtable
endprimitive

primitive OR6M12RA_udp_0(Z,A, B, C, D, E, F);
  output Z;
  input A, B, C, D, E, F;
  table
  //A, B, C, D, E, F: Z
    1  ?  ?  ?  ?  ?: 1;
    ?  1  ?  ?  ?  ?: 1;
    ?  ?  1  ?  ?  ?: 1;
    ?  ?  ?  1  ?  ?: 1;
    ?  ?  ?  ?  1  ?: 1;
    ?  ?  ?  ?  ?  1: 1;
    0  0  0  0  0  0: 0;
  endtable
endprimitive

primitive REG1M1R_udp_0(MGM_WB_0,IQN, RG, RGB);
  output MGM_WB_0;
  input IQN, RG, RGB;
  table
  //IQN, RG, RGB: MGM_WB_0
    1  1  0: 1;
    0  1  0: 0;
    ?  0  0: 1;
    ?  0  1: 1;
    ?  1  1: 1;
  endtable
endprimitive

primitive SDFAQM1RA_udp_0(MGM_D,A, B, SE, SD);
  output MGM_D;
  input A, B, SE, SD;
  table
  //A, B, SE, SD: MGM_D
    1  1  0  ?: 1;
    ?  ?  1  1: 1;
    0  ?  0  ?: 0;
    ?  0  0  ?: 0;
    ?  ?  1  0: 0;
    1  1  ?  1: 1;
    0  ?  ?  0: 0;
    ?  0  ?  0: 0;
  endtable
endprimitive

primitive SDFEM1RA_udp_0(MGM_D,D, E, SE, IQ, SD);
  output MGM_D;
  input D, E, SE, IQ, SD;
  table
  //D, E, SE, IQ, SD: MGM_D
    1  1  0  ?  ?: 1;
    1  ?  0  1  ?: 1;
    ?  0  0  1  ?: 1;
    ?  ?  1  ?  1: 1;
    0  1  0  ?  ?: 0;
    0  ?  0  0  ?: 0;
    ?  0  0  0  ?: 0;
    ?  ?  1  ?  0: 0;
    1  1  ?  ?  1: 1;
    1  ?  ?  1  1: 1;
    ?  0  ?  1  1: 1;
    0  1  ?  ?  0: 0;
    0  ?  ?  0  0: 0;
    ?  0  ?  0  0: 0;
  endtable
endprimitive

primitive SDFEQZRM1RA_udp_0(MGM_D,D, E, RB, SE, IQ, SD);
  output MGM_D;
  input D, E, RB, SE, IQ, SD;
  table
  //D, E, RB, SE, IQ, SD: MGM_D
    1  1  1  0  ?  ?: 1;
    1  ?  1  0  1  ?: 1;
    ?  0  1  0  1  ?: 1;
    ?  ?  ?  1  ?  1: 1;
    0  1  ?  0  ?  ?: 0;
    0  ?  ?  0  0  ?: 0;
    ?  0  ?  0  0  ?: 0;
    ?  ?  0  0  ?  ?: 0;
    ?  ?  ?  1  ?  0: 0;
    1  1  1  ?  ?  1: 1;
    1  ?  1  ?  1  1: 1;
    ?  0  1  ?  1  1: 1;
    0  1  ?  ?  ?  0: 0;
    0  ?  ?  ?  0  0: 0;
    ?  0  ?  ?  0  0: 0;
    ?  ?  0  ?  ?  0: 0;
  endtable
endprimitive

primitive SDFMM1RA_udp_0(MGM_D,D1, S, SE, D2, SD);
  output MGM_D;
  input D1, S, SE, D2, SD;
  table
  //D1, S, SE, D2, SD: MGM_D
    1  1  0  ?  ?: 1;
    ?  0  0  1  ?: 1;
    ?  ?  1  ?  1: 1;
    0  1  0  ?  ?: 0;
    ?  0  0  0  ?: 0;
    ?  ?  1  ?  0: 0;
    1  1  ?  ?  1: 1;
    ?  0  ?  1  1: 1;
    0  1  ?  ?  0: 0;
    ?  0  ?  0  0: 0;
    1  ?  0  1  ?: 1;
    0  ?  0  0  ?: 0;
    1  ?  ?  1  1: 1;
    0  ?  ?  0  0: 0;
  endtable
endprimitive

primitive SDFQZRSM1RA_udp_0(MGM_D,D, RB, SE, SB, SD);
  output MGM_D;
  input D, RB, SE, SB, SD;
  table
  //D, RB, SE, SB, SD: MGM_D
    1  1  0  ?  ?: 1;
    ?  1  0  0  ?: 1;
    ?  ?  1  ?  1: 1;
    0  ?  0  1  ?: 0;
    ?  0  0  ?  ?: 0;
    ?  ?  1  ?  0: 0;
    1  1  ?  ?  1: 1;
    ?  1  ?  0  1: 1;
    0  ?  ?  1  0: 0;
    ?  0  ?  ?  0: 0;
  endtable
endprimitive

primitive SDFQZSM1RA_udp_0(MGM_D,D, SE, SB, SD);
  output MGM_D;
  input D, SE, SB, SD;
  table
  //D, SE, SB, SD: MGM_D
    1  0  ?  ?: 1;
    ?  0  0  ?: 1;
    ?  1  ?  1: 1;
    0  0  1  ?: 0;
    ?  1  ?  0: 0;
    1  ?  ?  1: 1;
    ?  ?  0  1: 1;
    0  ?  1  0: 0;
  endtable
endprimitive

primitive XNR4M1RA_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  1  1  1: 1;
    1  1  0  0: 1;
    1  0  1  0: 1;
    1  0  0  1: 1;
    0  1  1  0: 1;
    0  1  0  1: 1;
    0  0  1  1: 1;
    0  0  0  0: 1;
    1  1  1  0: 0;
    1  1  0  1: 0;
    1  0  1  1: 0;
    1  0  0  0: 0;
    0  1  1  1: 0;
    0  1  0  0: 0;
    0  0  1  0: 0;
    0  0  0  1: 0;
  endtable
endprimitive

primitive XOR4M1RA_udp_0(Z,A, B, C, D);
  output Z;
  input A, B, C, D;
  table
  //A, B, C, D: Z
    1  1  1  0: 1;
    1  1  0  1: 1;
    1  0  1  1: 1;
    1  0  0  0: 1;
    0  1  1  1: 1;
    0  1  0  0: 1;
    0  0  1  0: 1;
    0  0  0  1: 1;
    1  1  1  1: 0;
    1  1  0  0: 0;
    1  0  1  0: 0;
    1  0  0  1: 0;
    0  1  1  0: 0;
    0  1  0  1: 0;
    0  0  1  1: 0;
    0  0  0  0: 0;
  endtable
endprimitive
