--!
--! @file fll_top.vhd
--! @brief Frequency Locked Loop Top Level 
--! 
--! This is the top level of the Frequency Locked Loop (FLL)
--! This integrates the control part, the DCO, the clock counter, and the clock divider
--! 
--! <B>
--! @n
--! This file is part of the Platform 2012 program,
--! a cooperation between STMicroelectronics and CEA.@n
--! Redistribution of this file to outside parties is
--! strictly prohibited without the written consent
--! of the module owner indicated below.@n
--! </B>
--! 
--! @par  Module owner: Ivan MIRO PANADES
--!       ivan.miro-panades@cea.fr
--! 
--! @par  Copyright (C) 2009 CEA
--! 
--! @par  Authors:  Ivan MIRO PANADES
--!                 Pascal VIVET
--! 
--! @par  Id: $Id: fll_top.vhd 1 2014-01-15 16:11:08Z im219746 $
--! @par  Date: $Date: 2014-01-15 17:11:08 +0100 (Wed, 15 Jan 2014) $
--! @par  Revision: $Rev: 1 $
--!


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY common_cells_lib;
USE common_cells_lib.ALL;

ENTITY fll_top IS
  GENERIC (
    BYPASS_CMD_AFTER_RESET : STD_LOGIC_VECTOR(7 downto 0) := "10000000";
    CLK_DIV_AFTER_RESET    : STD_LOGIC_VECTOR := "0101"  -- Value aplied to the muxes at reset 
  );
  PORT(
    -- General signals
    rst_n               : IN  STD_LOGIC;                    -- reset, already re-synchronized with the CVP clock : clk
    rst_ref_n           : IN  STD_LOGIC;                    -- reset, already re-synchronized with the clk_ref clock 
    rst_async_n         : IN  STD_LOGIC;                    -- hard reset, fully asynchronous (used by fll_counter and fll_clk_ref)
    clk                 : IN  STD_LOGIC;                    -- CVP clock (~ 1GHz)
    clk_ref             : IN  STD_LOGIC;                    -- external reference clock (= 100MHz)
    enable              : IN  STD_LOGIC;
    test_mode           : IN  STD_LOGIC;                    -- test_mode : only DFT on the control block (clk domain)
    test_se             : IN  STD_LOGIC;
    --test_si             : IN  STD_LOGIC;
    --test_so             : OUT STD_LOGIC;
    
    -- configuration values
    cfg_done            : IN  STD_LOGIC;                    -- a new configuration is done, update the loop control
    cfg_gain            : IN  STD_LOGIC_VECTOR(8 downto 0); -- gain value (unsigned 9bit, fixed point, 7 fraction bits, value from 0 to 3.99)
    cfg_set_point       : IN  STD_LOGIC_VECTOR(7 downto 0); -- set-point value (unsigned 8bit, from 0 to 255)
    cfg_sample_clocks   : IN  STD_LOGIC_VECTOR(3 downto 0); -- nb cycles the sampling is done (from 0 to 15, default is 5)
    cfg_capture_clocks  : IN  STD_LOGIC_VECTOR(3 downto 0); -- nb cycles the capture is done (from 0 to 15, default is 15)
    cfg_init            : IN  STD_LOGIC;                    -- a new init is done, re-init the loop control 
    cfg_init_command    : IN  STD_LOGIC_VECTOR(7 downto 0); -- init command for freq to DCO (unsigned 8bit, from 0 to 255)
    cfg_nb_multi_cycles : IN  STD_LOGIC_VECTOR(2 downto 0); -- number of multi-cycles path for combinational logic (1..7 range, default is 4)
    cfg_bypass          : IN  STD_LOGIC;                    -- bypass control signal
    cfg_bypass_command  : IN  STD_LOGIC_VECTOR(7 downto 0); -- bypass command for direct DCO control (unsigned 8bit, from 0 to 255)
    cfg_div             : IN  STD_LOGIC_VECTOR(3 downto 0); -- config to select the DCO division factor (2^0 to 2^15)

    -- outputs
    measure_value       : OUT STD_LOGIC_VECTOR(7 downto 0); -- measure value (unsigned 8bit, from 0 to 255)
    error_value         : OUT STD_LOGIC_VECTOR(8 downto 0); -- error value (signed 9bit, from -256 to 255)
    dco_value           : OUT STD_LOGIC_VECTOR(7 downto 0); -- DCO applied value (unsigned 8bit, from 0 to 255)
    valid_clk           : OUT STD_LOGIC;                    -- output control to indicate that generated clock is now stable
    new_value_to_dco    : OUT STD_LOGIC;                    -- Generate a pulse on each new value to DCO
    current_set_point   : OUT STD_LOGIC_VECTOR(7 downto 0); -- current set_point
    current_div         : OUT STD_LOGIC_VECTOR(3 downto 0); -- current division factor
    clk_out             : OUT STD_LOGIC                     -- generated clock
  );
END fll_top;


ARCHITECTURE rtl of fll_top IS 

  ----------------------------------------------------------------------
  -- Signals/contants declarations -------------------------------------
  ----------------------------------------------------------------------

  SIGNAL clk_dco, clk_dco_i : STD_LOGIC;                    -- clock generated by the DCO

  SIGNAL freq_to_dco        : STD_LOGIC_VECTOR(7 downto 0); -- control to DCO (unsigned 8bit, from 0 to 255)
  SIGNAL counter            : STD_LOGIC_VECTOR(7 downto 0); -- counter value from DCO (unsigned 8bit, from 0 to 255)

  SIGNAL sample_ref         : STD_LOGIC;                    -- control signals to the FLL sampleer
  SIGNAL sample_counter     : STD_LOGIC;
  SIGNAL clear              : STD_LOGIC;

  SIGNAL clk_out_s          : STD_LOGIC;
  SIGNAL clk_out_buf        : STD_LOGIC;

  SIGNAL clk_cg_dco         : STD_LOGIC;
  SIGNAL enable_cg_dco      : STD_LOGIC;
  SIGNAL new_value_to_dco_i : STD_LOGIC;

  SIGNAL enable_with_reset  : STD_LOGIC;
  
  ----------------------------------------------------------------------
  -- Components declarations -------------------------------------------
  ----------------------------------------------------------------------

  COMPONENT fll_clk_ref IS
    PORT(
      rst_ref_n      : IN  STD_LOGIC;                    -- hard reset
      clk_ref        : IN  STD_LOGIC;                    -- external reference clock (= 100MHz)
      test_mode      : IN  STD_LOGIC;                    -- test_mode from CVP
      sample_clocks  : IN  STD_LOGIC_VECTOR(3 downto 0); -- nb cycles the sampling is done (from 0 to 15, default is 5)
      capture_clocks : IN  STD_LOGIC_VECTOR(3 downto 0); -- nb cycles the capture is done (from 0 to 15, default is 15)
      sample         : OUT STD_LOGIC                     -- sample signal to clock counter
    );
  END COMPONENT;

  COMPONENT fll_control IS
    GENERIC (
      BYPASS_CMD_AFTER_RESET : STD_LOGIC_VECTOR(7 downto 0) := "10000000"
    );
    PORT(
      -- General signals
      rst_n             : IN  STD_LOGIC;
      clk               : IN  STD_LOGIC;                      -- this is the CVP clock (~ 1GHz)
      test_mode         : IN  STD_LOGIC;                      -- test_mode from CVP
  
      -- configuration values
      cfg_done          : IN  STD_LOGIC;                      -- a new configuration is done, update the loop control 
      cfg_gain          : IN  STD_LOGIC_VECTOR(8 downto 0);   -- gain value (unsigned 9bit, fixed point, 7 fraction bits, value from 0 to 3.99)
      cfg_set_point     : IN  STD_LOGIC_VECTOR(7 downto 0);   -- set-point value (unsigned 8bit, from 0 to 255)
      cfg_init          : IN  STD_LOGIC;                      -- a new init is done, re-init the loop control
      cfg_init_command  : IN  STD_LOGIC_VECTOR(7 downto 0);   -- init command for freq to DCO (unsigned 8bit, from 0 to 255)
      cfg_nb_multi_cycles : IN  STD_LOGIC_VECTOR(2 downto 0); -- number of multi-cycles path for combinational logic (2..7 range, default is 4)
      cfg_bypass        : IN  STD_LOGIC;                      -- bypass control signal
      cfg_bypass_command: IN  STD_LOGIC_VECTOR(7 downto 0);   -- bypass command for direct DCO control (unsigned 8bit, from 0 to 255)
  
      -- From/To counter module
      sample            : IN  STD_LOGIC;                      -- sample signal from counter
      counter           : IN  STD_LOGIC_VECTOR(7 downto 0);   -- counter value from DCO (unsigned 8bit, from 0 to 255)
      clear             : OUT STD_LOGIC;                      -- clear signal back to the counter
  
      -- outputs
      new_value_to_dco  : OUT STD_LOGIC;                      -- Generate a pulse on each new value to DCO
      current_set_point : OUT STD_LOGIC_VECTOR(7 downto 0);   -- current set_point
      freq_to_dco       : OUT STD_LOGIC_VECTOR(7 downto 0);   -- control to DCO (unsigned 8bit, from 0 to 255)
      dco_value         : OUT STD_LOGIC_VECTOR(7 downto 0);   -- Current DCO value (unsigned 8bit, from 0 to 255)
      measure_value     : OUT STD_LOGIC_VECTOR(7 downto 0);   -- measure value (unsigned 8bit, from 0 to 255)
      error_value       : OUT STD_LOGIC_VECTOR(8 downto 0)    -- error value (signed 9bit, from -256 to 255)
    );
  END COMPONENT;

  COMPONENT DCO IS
    PORT(
      FREQ   : IN  STD_LOGIC_VECTOR(7 downto 0);
      TI     : IN  STD_LOGIC;
      TE     : IN  STD_LOGIC;
      CP     : IN  STD_LOGIC;
      RN     : IN  STD_LOGIC;
      ENAB   : IN  STD_LOGIC;
      TQ     : OUT STD_LOGIC;
      FOUT   : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT fll_counter IS
    PORT(
      clk_dco        : IN  STD_LOGIC;                    -- clk generated by VCO/DCO
      rst_async_n    : IN  STD_LOGIC;                    -- hard reset
      test_mode      : IN  STD_LOGIC;                    -- test_mode from CVP
      clear          : IN  STD_LOGIC;                    -- clear input signal
      sample_i       : IN  STD_LOGIC;                    -- sample input signal, set during NB cycles clk_ref
      sample_o       : OUT STD_LOGIC;                    -- sample output signal, resynchronized with clk_dco
      counter        : OUT STD_LOGIC_VECTOR(7 downto 0)  -- counter value, send back to control
    );
  END COMPONENT;

  COMPONENT fll_clk_div_select IS
    GENERIC(
      CLK_DIV_AFTER_RESET : STD_LOGIC_VECTOR := "1000"  -- Value aplied to the muxes at reset 
    );
    PORT(
      clk          : IN  STD_LOGIC;                    -- Main clock (CVP)
      clk_dco      : IN  STD_LOGIC;                    -- clk generated by the VCO/DCO
      rst_n        : IN  STD_LOGIC;                    -- reset already synchronized within CVP
      rst_async_n  : IN  STD_LOGIC;                    -- hard reset
      cfg_div      : IN  STD_LOGIC_VECTOR(3 downto 0); -- config to select the DCO division factor (2^0 to 2^15)
      test_mode    : IN  STD_LOGIC;
      clk_out      : OUT STD_LOGIC;                    -- generated clock
      valid_clk    : OUT STD_LOGIC;                    -- output control to indicate that generated clock is now stable
      current_div  : OUT STD_LOGIC_VECTOR(3 downto 0)  -- current division factor
      ); 
  END COMPONENT;
    
  COMPONENT clock_mux2 IS
    PORT(
      clk_in0     : IN  STD_LOGIC;
      clk_in1     : IN  STD_LOGIC;
      clk_select  : IN  STD_LOGIC;
      clk_out     : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT clock_buffer IS
    PORT(
      clk_in      : IN  STD_LOGIC;
      clk_out     : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT clock_gating IS
    PORT(
      clk_in      : IN  STD_LOGIC;
      enable      : IN  STD_LOGIC;
      test_mode   : IN  STD_LOGIC;
      clk_out     : OUT STD_LOGIC
    );
  END COMPONENT;


BEGIN

  --------------------------------------------------------------------------------
  -- FLL clk ref
  --------------------------------------------------------------------------------

  fll_clk_ref_u : fll_clk_ref 
    PORT MAP (
        rst_ref_n      => rst_ref_n ,       
        clk_ref        => clk_ref,  -- external reference clock (= 100MHz)
        test_mode      => test_mode     ,
        sample_clocks  => cfg_sample_clocks ,
        capture_clocks => cfg_capture_clocks,
        sample         => sample_ref       -- sample signal to clock counter
    );

  --------------------------------------------------------------------------------
  -- FLL Control
  --------------------------------------------------------------------------------

  fll_control_u : fll_control
    GENERIC MAP (
      BYPASS_CMD_AFTER_RESET => BYPASS_CMD_AFTER_RESET
    )
    PORT MAP (
      -- General signals
      rst_n               => rst_n  ,
      clk                 => clk      ,
      test_mode           => test_mode,

      -- configuration values
      cfg_done            => cfg_done           ,
      cfg_gain            => cfg_gain           ,
      cfg_set_point       => cfg_set_point      ,
      cfg_init            => cfg_init           ,
      cfg_init_command    => cfg_init_command   ,
      cfg_nb_multi_cycles => cfg_nb_multi_cycles,
      cfg_bypass          => cfg_bypass         ,
      cfg_bypass_command  => cfg_bypass_command ,

      -- From/To counter module
      sample              => sample_counter,         
      counter             => counter       ,
      clear               => clear         ,
    
      -- outputs        -- outputs
      new_value_to_dco    => new_value_to_dco_i,
      current_set_point   => current_set_point,
      freq_to_dco         => freq_to_dco  ,      
      dco_value           => dco_value,
      measure_value       => measure_value,
      error_value         => error_value  
      );


  --------------------------------------------------------------------------------
  -- FLL DCO
  --------------------------------------------------------------------------------
  u_cg_DCO : clock_gating
    PORT MAP(
      clk_in     => clk,
      enable     => enable_cg_dco,
      test_mode  => test_mode,
      clk_out    => clk_cg_dco
    );

  enable_cg_dco <= new_value_to_dco_i OR cfg_bypass;

  fll_dco_u : DCO
    PORT MAP (
      FREQ  => freq_to_dco,
      TI    => '0', 
      TE    => test_se, 
      CP    => clk_cg_dco,
      RN    => rst_n, 
      ENAB  => enable_with_reset,
      TQ    => open, 
      FOUT  => clk_dco
    );
  
  --When reset is active, the DCO is also in reset
  enable_with_reset <= enable AND rst_async_n;

  --------------------------------------------------------------------------------
  -- Clock mux for testability
  --------------------------------------------------------------------------------
  clk_mux_for_test_u : clock_mux2 
    PORT MAP(
      clk_in0     => clk_dco  ,
      clk_in1     => clk      ,
      clk_select  => test_mode,
      clk_out     => clk_dco_i
    );

  --------------------------------------------------------------------------------
  -- FLL Counter
  --------------------------------------------------------------------------------

  fll_counter_u : fll_counter
    PORT MAP (
      clk_dco        => clk_dco_i , -- clk generated by VCO/DCO
      rst_async_n    => rst_async_n , -- hard reset
      test_mode      => test_mode     ,
      clear          => clear         ,
      sample_i       => sample_ref    , -- update=1 during 6th clk_ref
      sample_o       => sample_counter, -- update signal, resynchronized with clk_dco
      counter        => counter         -- counter value, send back to control
    );


  --------------------------------------------------------------------------------
  -- FLL clock divider and selector
  --------------------------------------------------------------------------------

  fll_clk_div_select_u : fll_clk_div_select
    GENERIC MAP(
      CLK_DIV_AFTER_RESET => CLK_DIV_AFTER_RESET  -- Value aplied to the muxes at reset 
    )
    PORT MAP(
      clk         => clk, 
      clk_dco     => clk_dco_i, 
      rst_n       => rst_n, 
      rst_async_n => rst_async_n, 
      cfg_div     => cfg_div, 
      test_mode   => test_mode, 
      clk_out     => clk_out_s, 
      valid_clk   => valid_clk,
      current_div => current_div
      );

  -- Clock buffer to break the timing loops if FLL output clock is used as FLL main clock 
  clk_buf_u : clock_buffer
    PORT MAP(
      clk_in    => clk_out_s,  
      clk_out   => clk_out_buf  
    );
  
  --Outputs
  clk_out   <= clk_out_buf;
  new_value_to_dco <= new_value_to_dco_i;
  
END rtl;

