module vbbgen_PULPV3_weakdriver
(
	input logic 		selP0,
	input logic 		selP1,
	input logic 		selN0,
	input logic 		selN1,
	input logic 		clk
);

endmodule // driverCombined
