`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO112X17_A_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X17_A_F_Z_F_100 0.1
`define C12T32_LLUP0_AO112X17_B_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X17_B_F_Z_F_100 0.1
`define C12T32_LLUP0_AO112X17_C_R_Z_R_010 0.1
`define C12T32_LLUP0_AO112X17_C_F_Z_F_010 0.1
`define C12T32_LLUP0_AO112X17_C_R_Z_R_000 0.1
`define C12T32_LLUP0_AO112X17_C_F_Z_F_000 0.1
`define C12T32_LLUP0_AO112X17_C_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X17_C_F_Z_F_100 0.1
`define C12T32_LLUP0_AO112X17_D_R_Z_R_010 0.1
`define C12T32_LLUP0_AO112X17_D_F_Z_F_010 0.1
`define C12T32_LLUP0_AO112X17_D_R_Z_R_000 0.1
`define C12T32_LLUP0_AO112X17_D_F_Z_F_000 0.1
`define C12T32_LLUP0_AO112X17_D_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X17_D_F_Z_F_100 0.1

module C12T32_LLUP0_AO112X17 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	and    U1 (INTERNAL1, A, B) ;
	or   #1 U2 (Z, INTERNAL1, C, D) ;



	specify

		if (B && !C && !D) (A +=> Z) = (`C12T32_LLUP0_AO112X17_A_R_Z_R_100,`C12T32_LLUP0_AO112X17_A_F_Z_F_100);
		if (A && !C && !D) (B +=> Z) = (`C12T32_LLUP0_AO112X17_B_R_Z_R_100,`C12T32_LLUP0_AO112X17_B_F_Z_F_100);
		if (!A && B && !D) (C +=> Z) = (`C12T32_LLUP0_AO112X17_C_R_Z_R_010,`C12T32_LLUP0_AO112X17_C_F_Z_F_010);
		if (!A && !B && !D) (C +=> Z) = (`C12T32_LLUP0_AO112X17_C_R_Z_R_000,`C12T32_LLUP0_AO112X17_C_F_Z_F_000);
		if (A && !B && !D) (C +=> Z) = (`C12T32_LLUP0_AO112X17_C_R_Z_R_100,`C12T32_LLUP0_AO112X17_C_F_Z_F_100);
		if (!A && B && !C) (D +=> Z) = (`C12T32_LLUP0_AO112X17_D_R_Z_R_010,`C12T32_LLUP0_AO112X17_D_F_Z_F_010);
		if (!A && !B && !C) (D +=> Z) = (`C12T32_LLUP0_AO112X17_D_R_Z_R_000,`C12T32_LLUP0_AO112X17_D_F_Z_F_000);
		if (A && !B && !C) (D +=> Z) = (`C12T32_LLUP0_AO112X17_D_R_Z_R_100,`C12T32_LLUP0_AO112X17_D_F_Z_F_100);


	endspecify

endmodule // C12T32_LLUP0_AO112X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO112X8_A_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X8_A_F_Z_F_100 0.1
`define C12T32_LLUP0_AO112X8_B_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X8_B_F_Z_F_100 0.1
`define C12T32_LLUP0_AO112X8_C_R_Z_R_010 0.1
`define C12T32_LLUP0_AO112X8_C_F_Z_F_010 0.1
`define C12T32_LLUP0_AO112X8_C_R_Z_R_000 0.1
`define C12T32_LLUP0_AO112X8_C_F_Z_F_000 0.1
`define C12T32_LLUP0_AO112X8_C_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X8_C_F_Z_F_100 0.1
`define C12T32_LLUP0_AO112X8_D_R_Z_R_010 0.1
`define C12T32_LLUP0_AO112X8_D_F_Z_F_010 0.1
`define C12T32_LLUP0_AO112X8_D_R_Z_R_000 0.1
`define C12T32_LLUP0_AO112X8_D_F_Z_F_000 0.1
`define C12T32_LLUP0_AO112X8_D_R_Z_R_100 0.1
`define C12T32_LLUP0_AO112X8_D_F_Z_F_100 0.1

module C12T32_LLUP0_AO112X8 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	and    U1 (INTERNAL1, A, B) ;
	or   #1 U2 (Z, INTERNAL1, C, D) ;



	specify

		if (B && !C && !D) (A +=> Z) = (`C12T32_LLUP0_AO112X8_A_R_Z_R_100,`C12T32_LLUP0_AO112X8_A_F_Z_F_100);
		if (A && !C && !D) (B +=> Z) = (`C12T32_LLUP0_AO112X8_B_R_Z_R_100,`C12T32_LLUP0_AO112X8_B_F_Z_F_100);
		if (!A && B && !D) (C +=> Z) = (`C12T32_LLUP0_AO112X8_C_R_Z_R_010,`C12T32_LLUP0_AO112X8_C_F_Z_F_010);
		if (!A && !B && !D) (C +=> Z) = (`C12T32_LLUP0_AO112X8_C_R_Z_R_000,`C12T32_LLUP0_AO112X8_C_F_Z_F_000);
		if (A && !B && !D) (C +=> Z) = (`C12T32_LLUP0_AO112X8_C_R_Z_R_100,`C12T32_LLUP0_AO112X8_C_F_Z_F_100);
		if (!A && B && !C) (D +=> Z) = (`C12T32_LLUP0_AO112X8_D_R_Z_R_010,`C12T32_LLUP0_AO112X8_D_F_Z_F_010);
		if (!A && !B && !C) (D +=> Z) = (`C12T32_LLUP0_AO112X8_D_R_Z_R_000,`C12T32_LLUP0_AO112X8_D_F_Z_F_000);
		if (A && !B && !C) (D +=> Z) = (`C12T32_LLUP0_AO112X8_D_R_Z_R_100,`C12T32_LLUP0_AO112X8_D_F_Z_F_100);


	endspecify

endmodule // C12T32_LLUP0_AO112X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO12X17_A_R_Z_R_10 0.1
`define C12T32_LLUP0_AO12X17_A_F_Z_F_10 0.1
`define C12T32_LLUP0_AO12X17_B_R_Z_R_10 0.1
`define C12T32_LLUP0_AO12X17_B_F_Z_F_10 0.1
`define C12T32_LLUP0_AO12X17_C_R_Z_R_00 0.1
`define C12T32_LLUP0_AO12X17_C_F_Z_F_00 0.1
`define C12T32_LLUP0_AO12X17_C_R_Z_R_10 0.1
`define C12T32_LLUP0_AO12X17_C_F_Z_F_10 0.1
`define C12T32_LLUP0_AO12X17_C_R_Z_R_01 0.1
`define C12T32_LLUP0_AO12X17_C_F_Z_F_01 0.1

module C12T32_LLUP0_AO12X17 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B) ;
	or   #1 U2 (Z, INTERNAL1, C) ;



	specify

		if (B && !C) (A +=> Z) = (`C12T32_LLUP0_AO12X17_A_R_Z_R_10,`C12T32_LLUP0_AO12X17_A_F_Z_F_10);
		if (A && !C) (B +=> Z) = (`C12T32_LLUP0_AO12X17_B_R_Z_R_10,`C12T32_LLUP0_AO12X17_B_F_Z_F_10);
		if (!A && !B) (C +=> Z) = (`C12T32_LLUP0_AO12X17_C_R_Z_R_00,`C12T32_LLUP0_AO12X17_C_F_Z_F_00);
		if (A && !B) (C +=> Z) = (`C12T32_LLUP0_AO12X17_C_R_Z_R_10,`C12T32_LLUP0_AO12X17_C_F_Z_F_10);
		if (!A && B) (C +=> Z) = (`C12T32_LLUP0_AO12X17_C_R_Z_R_01,`C12T32_LLUP0_AO12X17_C_F_Z_F_01);


	endspecify

endmodule // C12T32_LLUP0_AO12X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO12X8_A_R_Z_R_10 0.1
`define C12T32_LLUP0_AO12X8_A_F_Z_F_10 0.1
`define C12T32_LLUP0_AO12X8_B_R_Z_R_10 0.1
`define C12T32_LLUP0_AO12X8_B_F_Z_F_10 0.1
`define C12T32_LLUP0_AO12X8_C_R_Z_R_00 0.1
`define C12T32_LLUP0_AO12X8_C_F_Z_F_00 0.1
`define C12T32_LLUP0_AO12X8_C_R_Z_R_10 0.1
`define C12T32_LLUP0_AO12X8_C_F_Z_F_10 0.1
`define C12T32_LLUP0_AO12X8_C_R_Z_R_01 0.1
`define C12T32_LLUP0_AO12X8_C_F_Z_F_01 0.1

module C12T32_LLUP0_AO12X8 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B) ;
	or   #1 U2 (Z, INTERNAL1, C) ;



	specify

		if (B && !C) (A +=> Z) = (`C12T32_LLUP0_AO12X8_A_R_Z_R_10,`C12T32_LLUP0_AO12X8_A_F_Z_F_10);
		if (A && !C) (B +=> Z) = (`C12T32_LLUP0_AO12X8_B_R_Z_R_10,`C12T32_LLUP0_AO12X8_B_F_Z_F_10);
		if (!A && !B) (C +=> Z) = (`C12T32_LLUP0_AO12X8_C_R_Z_R_00,`C12T32_LLUP0_AO12X8_C_F_Z_F_00);
		if (A && !B) (C +=> Z) = (`C12T32_LLUP0_AO12X8_C_R_Z_R_10,`C12T32_LLUP0_AO12X8_C_F_Z_F_10);
		if (!A && B) (C +=> Z) = (`C12T32_LLUP0_AO12X8_C_R_Z_R_01,`C12T32_LLUP0_AO12X8_C_F_Z_F_01);


	endspecify

endmodule // C12T32_LLUP0_AO12X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO222X17_A_R_Z_R_11001 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_11001 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_11010 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_11010 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_11000 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_11000 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_10000 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_10000 0.1
`define C12T32_LLUP0_AO222X17_A_R_Z_R_10010 0.1
`define C12T32_LLUP0_AO222X17_A_F_Z_F_10010 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_11001 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_11001 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_11010 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_11010 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_11000 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_11000 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_10000 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_10000 0.1
`define C12T32_LLUP0_AO222X17_B_R_Z_R_10010 0.1
`define C12T32_LLUP0_AO222X17_B_F_Z_F_10010 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_01100 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_01100 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_01110 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_01110 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_00101 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_00100 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_00100 0.1
`define C12T32_LLUP0_AO222X17_C_R_Z_R_00110 0.1
`define C12T32_LLUP0_AO222X17_C_F_Z_F_00110 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_01100 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_01100 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_01110 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_01110 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_00101 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_00100 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_00100 0.1
`define C12T32_LLUP0_AO222X17_D_R_Z_R_00110 0.1
`define C12T32_LLUP0_AO222X17_D_F_Z_F_00110 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_10011 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_10011 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_01001 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_01001 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_01011 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_01011 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_00011 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_00011 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_00001 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_00001 0.1
`define C12T32_LLUP0_AO222X17_E_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X17_E_F_Z_F_00101 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_10011 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_10011 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_01001 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_01001 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_01011 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_01011 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_00011 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_00011 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_00001 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_00001 0.1
`define C12T32_LLUP0_AO222X17_F_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X17_F_F_Z_F_00101 0.1

module C12T32_LLUP0_AO222X17 (Z, A, B, C, D, E, F);

	output Z;
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;

	and    U1 (INTERNAL1, A, B) ;
	and    U2 (INTERNAL2, C, D) ;
	and    U3 (INTERNAL3, E, F) ;
	or   #1 U4 (Z, INTERNAL1, INTERNAL2, INTERNAL3) ;



	specify

		if (B && C && !D && !E && F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_11001,`C12T32_LLUP0_AO222X17_A_F_Z_F_11001);
		if (B && C && !D && E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_11010,`C12T32_LLUP0_AO222X17_A_F_Z_F_11010);
		if (B && !C && D && !E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_10100,`C12T32_LLUP0_AO222X17_A_F_Z_F_10100);
		if (B && !C && D && E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_10110,`C12T32_LLUP0_AO222X17_A_F_Z_F_10110);
		if (B && !C && D && !E && F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_10101,`C12T32_LLUP0_AO222X17_A_F_Z_F_10101);
		if (B && C && !D && !E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_11000,`C12T32_LLUP0_AO222X17_A_F_Z_F_11000);
		if (B && !C && !D && !E && F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_10001,`C12T32_LLUP0_AO222X17_A_F_Z_F_10001);
		if (B && !C && !D && !E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_10000,`C12T32_LLUP0_AO222X17_A_F_Z_F_10000);
		if (B && !C && !D && E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X17_A_R_Z_R_10010,`C12T32_LLUP0_AO222X17_A_F_Z_F_10010);
		if (A && C && !D && !E && F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_11001,`C12T32_LLUP0_AO222X17_B_F_Z_F_11001);
		if (A && C && !D && E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_11010,`C12T32_LLUP0_AO222X17_B_F_Z_F_11010);
		if (A && !C && D && !E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_10100,`C12T32_LLUP0_AO222X17_B_F_Z_F_10100);
		if (A && !C && D && E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_10110,`C12T32_LLUP0_AO222X17_B_F_Z_F_10110);
		if (A && !C && D && !E && F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_10101,`C12T32_LLUP0_AO222X17_B_F_Z_F_10101);
		if (A && C && !D && !E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_11000,`C12T32_LLUP0_AO222X17_B_F_Z_F_11000);
		if (A && !C && !D && !E && F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_10001,`C12T32_LLUP0_AO222X17_B_F_Z_F_10001);
		if (A && !C && !D && !E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_10000,`C12T32_LLUP0_AO222X17_B_F_Z_F_10000);
		if (A && !C && !D && E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X17_B_R_Z_R_10010,`C12T32_LLUP0_AO222X17_B_F_Z_F_10010);
		if (A && !B && D && !E && F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_10101,`C12T32_LLUP0_AO222X17_C_F_Z_F_10101);
		if (A && !B && D && E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_10110,`C12T32_LLUP0_AO222X17_C_F_Z_F_10110);
		if (!A && B && D && !E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_01100,`C12T32_LLUP0_AO222X17_C_F_Z_F_01100);
		if (!A && B && D && E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_01110,`C12T32_LLUP0_AO222X17_C_F_Z_F_01110);
		if (!A && B && D && !E && F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_01101,`C12T32_LLUP0_AO222X17_C_F_Z_F_01101);
		if (A && !B && D && !E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_10100,`C12T32_LLUP0_AO222X17_C_F_Z_F_10100);
		if (!A && !B && D && !E && F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_00101,`C12T32_LLUP0_AO222X17_C_F_Z_F_00101);
		if (!A && !B && D && !E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_00100,`C12T32_LLUP0_AO222X17_C_F_Z_F_00100);
		if (!A && !B && D && E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X17_C_R_Z_R_00110,`C12T32_LLUP0_AO222X17_C_F_Z_F_00110);
		if (A && !B && C && !E && F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_10101,`C12T32_LLUP0_AO222X17_D_F_Z_F_10101);
		if (A && !B && C && E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_10110,`C12T32_LLUP0_AO222X17_D_F_Z_F_10110);
		if (!A && B && C && !E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_01100,`C12T32_LLUP0_AO222X17_D_F_Z_F_01100);
		if (!A && B && C && E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_01110,`C12T32_LLUP0_AO222X17_D_F_Z_F_01110);
		if (!A && B && C && !E && F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_01101,`C12T32_LLUP0_AO222X17_D_F_Z_F_01101);
		if (A && !B && C && !E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_10100,`C12T32_LLUP0_AO222X17_D_F_Z_F_10100);
		if (!A && !B && C && !E && F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_00101,`C12T32_LLUP0_AO222X17_D_F_Z_F_00101);
		if (!A && !B && C && !E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_00100,`C12T32_LLUP0_AO222X17_D_F_Z_F_00100);
		if (!A && !B && C && E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X17_D_R_Z_R_00110,`C12T32_LLUP0_AO222X17_D_F_Z_F_00110);
		if (A && !B && !C && D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_10011,`C12T32_LLUP0_AO222X17_E_F_Z_F_10011);
		if (A && !B && C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_10101,`C12T32_LLUP0_AO222X17_E_F_Z_F_10101);
		if (!A && B && !C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_01001,`C12T32_LLUP0_AO222X17_E_F_Z_F_01001);
		if (!A && B && C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_01101,`C12T32_LLUP0_AO222X17_E_F_Z_F_01101);
		if (!A && B && !C && D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_01011,`C12T32_LLUP0_AO222X17_E_F_Z_F_01011);
		if (A && !B && !C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_10001,`C12T32_LLUP0_AO222X17_E_F_Z_F_10001);
		if (!A && !B && !C && D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_00011,`C12T32_LLUP0_AO222X17_E_F_Z_F_00011);
		if (!A && !B && !C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_00001,`C12T32_LLUP0_AO222X17_E_F_Z_F_00001);
		if (!A && !B && C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X17_E_R_Z_R_00101,`C12T32_LLUP0_AO222X17_E_F_Z_F_00101);
		if (A && !B && !C && D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_10011,`C12T32_LLUP0_AO222X17_F_F_Z_F_10011);
		if (A && !B && C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_10101,`C12T32_LLUP0_AO222X17_F_F_Z_F_10101);
		if (!A && B && !C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_01001,`C12T32_LLUP0_AO222X17_F_F_Z_F_01001);
		if (!A && B && C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_01101,`C12T32_LLUP0_AO222X17_F_F_Z_F_01101);
		if (!A && B && !C && D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_01011,`C12T32_LLUP0_AO222X17_F_F_Z_F_01011);
		if (A && !B && !C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_10001,`C12T32_LLUP0_AO222X17_F_F_Z_F_10001);
		if (!A && !B && !C && D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_00011,`C12T32_LLUP0_AO222X17_F_F_Z_F_00011);
		if (!A && !B && !C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_00001,`C12T32_LLUP0_AO222X17_F_F_Z_F_00001);
		if (!A && !B && C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X17_F_R_Z_R_00101,`C12T32_LLUP0_AO222X17_F_F_Z_F_00101);


	endspecify

endmodule // C12T32_LLUP0_AO222X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO222X8_A_R_Z_R_11001 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_11001 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_11010 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_11010 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_11000 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_11000 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_10000 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_10000 0.1
`define C12T32_LLUP0_AO222X8_A_R_Z_R_10010 0.1
`define C12T32_LLUP0_AO222X8_A_F_Z_F_10010 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_11001 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_11001 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_11010 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_11010 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_11000 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_11000 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_10000 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_10000 0.1
`define C12T32_LLUP0_AO222X8_B_R_Z_R_10010 0.1
`define C12T32_LLUP0_AO222X8_B_F_Z_F_10010 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_01100 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_01100 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_01110 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_01110 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_00101 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_00100 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_00100 0.1
`define C12T32_LLUP0_AO222X8_C_R_Z_R_00110 0.1
`define C12T32_LLUP0_AO222X8_C_F_Z_F_00110 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_10110 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_10110 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_01100 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_01100 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_01110 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_01110 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_10100 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_10100 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_00101 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_00100 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_00100 0.1
`define C12T32_LLUP0_AO222X8_D_R_Z_R_00110 0.1
`define C12T32_LLUP0_AO222X8_D_F_Z_F_00110 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_10011 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_10011 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_01001 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_01001 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_01011 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_01011 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_00011 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_00011 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_00001 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_00001 0.1
`define C12T32_LLUP0_AO222X8_E_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X8_E_F_Z_F_00101 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_10011 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_10011 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_10101 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_10101 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_01001 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_01001 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_01101 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_01101 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_01011 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_01011 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_10001 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_10001 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_00011 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_00011 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_00001 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_00001 0.1
`define C12T32_LLUP0_AO222X8_F_R_Z_R_00101 0.1
`define C12T32_LLUP0_AO222X8_F_F_Z_F_00101 0.1

module C12T32_LLUP0_AO222X8 (Z, A, B, C, D, E, F);

	output Z;
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;

	and    U1 (INTERNAL1, A, B) ;
	and    U2 (INTERNAL2, C, D) ;
	and    U3 (INTERNAL3, E, F) ;
	or   #1 U4 (Z, INTERNAL1, INTERNAL2, INTERNAL3) ;



	specify

		if (B && C && !D && !E && F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_11001,`C12T32_LLUP0_AO222X8_A_F_Z_F_11001);
		if (B && C && !D && E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_11010,`C12T32_LLUP0_AO222X8_A_F_Z_F_11010);
		if (B && !C && D && !E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_10100,`C12T32_LLUP0_AO222X8_A_F_Z_F_10100);
		if (B && !C && D && E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_10110,`C12T32_LLUP0_AO222X8_A_F_Z_F_10110);
		if (B && !C && D && !E && F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_10101,`C12T32_LLUP0_AO222X8_A_F_Z_F_10101);
		if (B && C && !D && !E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_11000,`C12T32_LLUP0_AO222X8_A_F_Z_F_11000);
		if (B && !C && !D && !E && F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_10001,`C12T32_LLUP0_AO222X8_A_F_Z_F_10001);
		if (B && !C && !D && !E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_10000,`C12T32_LLUP0_AO222X8_A_F_Z_F_10000);
		if (B && !C && !D && E && !F) (A +=> Z) = (`C12T32_LLUP0_AO222X8_A_R_Z_R_10010,`C12T32_LLUP0_AO222X8_A_F_Z_F_10010);
		if (A && C && !D && !E && F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_11001,`C12T32_LLUP0_AO222X8_B_F_Z_F_11001);
		if (A && C && !D && E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_11010,`C12T32_LLUP0_AO222X8_B_F_Z_F_11010);
		if (A && !C && D && !E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_10100,`C12T32_LLUP0_AO222X8_B_F_Z_F_10100);
		if (A && !C && D && E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_10110,`C12T32_LLUP0_AO222X8_B_F_Z_F_10110);
		if (A && !C && D && !E && F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_10101,`C12T32_LLUP0_AO222X8_B_F_Z_F_10101);
		if (A && C && !D && !E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_11000,`C12T32_LLUP0_AO222X8_B_F_Z_F_11000);
		if (A && !C && !D && !E && F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_10001,`C12T32_LLUP0_AO222X8_B_F_Z_F_10001);
		if (A && !C && !D && !E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_10000,`C12T32_LLUP0_AO222X8_B_F_Z_F_10000);
		if (A && !C && !D && E && !F) (B +=> Z) = (`C12T32_LLUP0_AO222X8_B_R_Z_R_10010,`C12T32_LLUP0_AO222X8_B_F_Z_F_10010);
		if (A && !B && D && !E && F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_10101,`C12T32_LLUP0_AO222X8_C_F_Z_F_10101);
		if (A && !B && D && E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_10110,`C12T32_LLUP0_AO222X8_C_F_Z_F_10110);
		if (!A && B && D && !E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_01100,`C12T32_LLUP0_AO222X8_C_F_Z_F_01100);
		if (!A && B && D && E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_01110,`C12T32_LLUP0_AO222X8_C_F_Z_F_01110);
		if (!A && B && D && !E && F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_01101,`C12T32_LLUP0_AO222X8_C_F_Z_F_01101);
		if (A && !B && D && !E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_10100,`C12T32_LLUP0_AO222X8_C_F_Z_F_10100);
		if (!A && !B && D && !E && F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_00101,`C12T32_LLUP0_AO222X8_C_F_Z_F_00101);
		if (!A && !B && D && !E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_00100,`C12T32_LLUP0_AO222X8_C_F_Z_F_00100);
		if (!A && !B && D && E && !F) (C +=> Z) = (`C12T32_LLUP0_AO222X8_C_R_Z_R_00110,`C12T32_LLUP0_AO222X8_C_F_Z_F_00110);
		if (A && !B && C && !E && F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_10101,`C12T32_LLUP0_AO222X8_D_F_Z_F_10101);
		if (A && !B && C && E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_10110,`C12T32_LLUP0_AO222X8_D_F_Z_F_10110);
		if (!A && B && C && !E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_01100,`C12T32_LLUP0_AO222X8_D_F_Z_F_01100);
		if (!A && B && C && E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_01110,`C12T32_LLUP0_AO222X8_D_F_Z_F_01110);
		if (!A && B && C && !E && F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_01101,`C12T32_LLUP0_AO222X8_D_F_Z_F_01101);
		if (A && !B && C && !E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_10100,`C12T32_LLUP0_AO222X8_D_F_Z_F_10100);
		if (!A && !B && C && !E && F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_00101,`C12T32_LLUP0_AO222X8_D_F_Z_F_00101);
		if (!A && !B && C && !E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_00100,`C12T32_LLUP0_AO222X8_D_F_Z_F_00100);
		if (!A && !B && C && E && !F) (D +=> Z) = (`C12T32_LLUP0_AO222X8_D_R_Z_R_00110,`C12T32_LLUP0_AO222X8_D_F_Z_F_00110);
		if (A && !B && !C && D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_10011,`C12T32_LLUP0_AO222X8_E_F_Z_F_10011);
		if (A && !B && C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_10101,`C12T32_LLUP0_AO222X8_E_F_Z_F_10101);
		if (!A && B && !C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_01001,`C12T32_LLUP0_AO222X8_E_F_Z_F_01001);
		if (!A && B && C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_01101,`C12T32_LLUP0_AO222X8_E_F_Z_F_01101);
		if (!A && B && !C && D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_01011,`C12T32_LLUP0_AO222X8_E_F_Z_F_01011);
		if (A && !B && !C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_10001,`C12T32_LLUP0_AO222X8_E_F_Z_F_10001);
		if (!A && !B && !C && D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_00011,`C12T32_LLUP0_AO222X8_E_F_Z_F_00011);
		if (!A && !B && !C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_00001,`C12T32_LLUP0_AO222X8_E_F_Z_F_00001);
		if (!A && !B && C && !D && F) (E +=> Z) = (`C12T32_LLUP0_AO222X8_E_R_Z_R_00101,`C12T32_LLUP0_AO222X8_E_F_Z_F_00101);
		if (A && !B && !C && D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_10011,`C12T32_LLUP0_AO222X8_F_F_Z_F_10011);
		if (A && !B && C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_10101,`C12T32_LLUP0_AO222X8_F_F_Z_F_10101);
		if (!A && B && !C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_01001,`C12T32_LLUP0_AO222X8_F_F_Z_F_01001);
		if (!A && B && C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_01101,`C12T32_LLUP0_AO222X8_F_F_Z_F_01101);
		if (!A && B && !C && D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_01011,`C12T32_LLUP0_AO222X8_F_F_Z_F_01011);
		if (A && !B && !C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_10001,`C12T32_LLUP0_AO222X8_F_F_Z_F_10001);
		if (!A && !B && !C && D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_00011,`C12T32_LLUP0_AO222X8_F_F_Z_F_00011);
		if (!A && !B && !C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_00001,`C12T32_LLUP0_AO222X8_F_F_Z_F_00001);
		if (!A && !B && C && !D && E) (F +=> Z) = (`C12T32_LLUP0_AO222X8_F_R_Z_R_00101,`C12T32_LLUP0_AO222X8_F_F_Z_F_00101);


	endspecify

endmodule // C12T32_LLUP0_AO222X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO22X17_A_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X17_A_F_Z_F_101 0.1
`define C12T32_LLUP0_AO22X17_A_R_Z_R_100 0.1
`define C12T32_LLUP0_AO22X17_A_F_Z_F_100 0.1
`define C12T32_LLUP0_AO22X17_A_R_Z_R_110 0.1
`define C12T32_LLUP0_AO22X17_A_F_Z_F_110 0.1
`define C12T32_LLUP0_AO22X17_B_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X17_B_F_Z_F_101 0.1
`define C12T32_LLUP0_AO22X17_B_R_Z_R_100 0.1
`define C12T32_LLUP0_AO22X17_B_F_Z_F_100 0.1
`define C12T32_LLUP0_AO22X17_B_R_Z_R_110 0.1
`define C12T32_LLUP0_AO22X17_B_F_Z_F_110 0.1
`define C12T32_LLUP0_AO22X17_C_R_Z_R_011 0.1
`define C12T32_LLUP0_AO22X17_C_F_Z_F_011 0.1
`define C12T32_LLUP0_AO22X17_C_R_Z_R_001 0.1
`define C12T32_LLUP0_AO22X17_C_F_Z_F_001 0.1
`define C12T32_LLUP0_AO22X17_C_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X17_C_F_Z_F_101 0.1
`define C12T32_LLUP0_AO22X17_D_R_Z_R_011 0.1
`define C12T32_LLUP0_AO22X17_D_F_Z_F_011 0.1
`define C12T32_LLUP0_AO22X17_D_R_Z_R_001 0.1
`define C12T32_LLUP0_AO22X17_D_F_Z_F_001 0.1
`define C12T32_LLUP0_AO22X17_D_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X17_D_F_Z_F_101 0.1

module C12T32_LLUP0_AO22X17 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	and    U1 (INTERNAL1, A, B) ;
	and    U2 (INTERNAL2, C, D) ;
	or   #1 U3 (Z, INTERNAL1, INTERNAL2) ;



	specify

		if (B && !C && D) (A +=> Z) = (`C12T32_LLUP0_AO22X17_A_R_Z_R_101,`C12T32_LLUP0_AO22X17_A_F_Z_F_101);
		if (B && !C && !D) (A +=> Z) = (`C12T32_LLUP0_AO22X17_A_R_Z_R_100,`C12T32_LLUP0_AO22X17_A_F_Z_F_100);
		if (B && C && !D) (A +=> Z) = (`C12T32_LLUP0_AO22X17_A_R_Z_R_110,`C12T32_LLUP0_AO22X17_A_F_Z_F_110);
		if (A && !C && D) (B +=> Z) = (`C12T32_LLUP0_AO22X17_B_R_Z_R_101,`C12T32_LLUP0_AO22X17_B_F_Z_F_101);
		if (A && !C && !D) (B +=> Z) = (`C12T32_LLUP0_AO22X17_B_R_Z_R_100,`C12T32_LLUP0_AO22X17_B_F_Z_F_100);
		if (A && C && !D) (B +=> Z) = (`C12T32_LLUP0_AO22X17_B_R_Z_R_110,`C12T32_LLUP0_AO22X17_B_F_Z_F_110);
		if (!A && B && D) (C +=> Z) = (`C12T32_LLUP0_AO22X17_C_R_Z_R_011,`C12T32_LLUP0_AO22X17_C_F_Z_F_011);
		if (!A && !B && D) (C +=> Z) = (`C12T32_LLUP0_AO22X17_C_R_Z_R_001,`C12T32_LLUP0_AO22X17_C_F_Z_F_001);
		if (A && !B && D) (C +=> Z) = (`C12T32_LLUP0_AO22X17_C_R_Z_R_101,`C12T32_LLUP0_AO22X17_C_F_Z_F_101);
		if (!A && B && C) (D +=> Z) = (`C12T32_LLUP0_AO22X17_D_R_Z_R_011,`C12T32_LLUP0_AO22X17_D_F_Z_F_011);
		if (!A && !B && C) (D +=> Z) = (`C12T32_LLUP0_AO22X17_D_R_Z_R_001,`C12T32_LLUP0_AO22X17_D_F_Z_F_001);
		if (A && !B && C) (D +=> Z) = (`C12T32_LLUP0_AO22X17_D_R_Z_R_101,`C12T32_LLUP0_AO22X17_D_F_Z_F_101);


	endspecify

endmodule // C12T32_LLUP0_AO22X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AO22X8_A_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X8_A_F_Z_F_101 0.1
`define C12T32_LLUP0_AO22X8_A_R_Z_R_100 0.1
`define C12T32_LLUP0_AO22X8_A_F_Z_F_100 0.1
`define C12T32_LLUP0_AO22X8_A_R_Z_R_110 0.1
`define C12T32_LLUP0_AO22X8_A_F_Z_F_110 0.1
`define C12T32_LLUP0_AO22X8_B_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X8_B_F_Z_F_101 0.1
`define C12T32_LLUP0_AO22X8_B_R_Z_R_100 0.1
`define C12T32_LLUP0_AO22X8_B_F_Z_F_100 0.1
`define C12T32_LLUP0_AO22X8_B_R_Z_R_110 0.1
`define C12T32_LLUP0_AO22X8_B_F_Z_F_110 0.1
`define C12T32_LLUP0_AO22X8_C_R_Z_R_011 0.1
`define C12T32_LLUP0_AO22X8_C_F_Z_F_011 0.1
`define C12T32_LLUP0_AO22X8_C_R_Z_R_001 0.1
`define C12T32_LLUP0_AO22X8_C_F_Z_F_001 0.1
`define C12T32_LLUP0_AO22X8_C_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X8_C_F_Z_F_101 0.1
`define C12T32_LLUP0_AO22X8_D_R_Z_R_011 0.1
`define C12T32_LLUP0_AO22X8_D_F_Z_F_011 0.1
`define C12T32_LLUP0_AO22X8_D_R_Z_R_001 0.1
`define C12T32_LLUP0_AO22X8_D_F_Z_F_001 0.1
`define C12T32_LLUP0_AO22X8_D_R_Z_R_101 0.1
`define C12T32_LLUP0_AO22X8_D_F_Z_F_101 0.1

module C12T32_LLUP0_AO22X8 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	and    U1 (INTERNAL1, A, B) ;
	and    U2 (INTERNAL2, C, D) ;
	or   #1 U3 (Z, INTERNAL1, INTERNAL2) ;



	specify

		if (B && !C && D) (A +=> Z) = (`C12T32_LLUP0_AO22X8_A_R_Z_R_101,`C12T32_LLUP0_AO22X8_A_F_Z_F_101);
		if (B && !C && !D) (A +=> Z) = (`C12T32_LLUP0_AO22X8_A_R_Z_R_100,`C12T32_LLUP0_AO22X8_A_F_Z_F_100);
		if (B && C && !D) (A +=> Z) = (`C12T32_LLUP0_AO22X8_A_R_Z_R_110,`C12T32_LLUP0_AO22X8_A_F_Z_F_110);
		if (A && !C && D) (B +=> Z) = (`C12T32_LLUP0_AO22X8_B_R_Z_R_101,`C12T32_LLUP0_AO22X8_B_F_Z_F_101);
		if (A && !C && !D) (B +=> Z) = (`C12T32_LLUP0_AO22X8_B_R_Z_R_100,`C12T32_LLUP0_AO22X8_B_F_Z_F_100);
		if (A && C && !D) (B +=> Z) = (`C12T32_LLUP0_AO22X8_B_R_Z_R_110,`C12T32_LLUP0_AO22X8_B_F_Z_F_110);
		if (!A && B && D) (C +=> Z) = (`C12T32_LLUP0_AO22X8_C_R_Z_R_011,`C12T32_LLUP0_AO22X8_C_F_Z_F_011);
		if (!A && !B && D) (C +=> Z) = (`C12T32_LLUP0_AO22X8_C_R_Z_R_001,`C12T32_LLUP0_AO22X8_C_F_Z_F_001);
		if (A && !B && D) (C +=> Z) = (`C12T32_LLUP0_AO22X8_C_R_Z_R_101,`C12T32_LLUP0_AO22X8_C_F_Z_F_101);
		if (!A && B && C) (D +=> Z) = (`C12T32_LLUP0_AO22X8_D_R_Z_R_011,`C12T32_LLUP0_AO22X8_D_F_Z_F_011);
		if (!A && !B && C) (D +=> Z) = (`C12T32_LLUP0_AO22X8_D_R_Z_R_001,`C12T32_LLUP0_AO22X8_D_F_Z_F_001);
		if (A && !B && C) (D +=> Z) = (`C12T32_LLUP0_AO22X8_D_R_Z_R_101,`C12T32_LLUP0_AO22X8_D_F_Z_F_101);


	endspecify

endmodule // C12T32_LLUP0_AO22X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_AOI21X11_A_R_Z_F_10 0.1
`define C12T32_LLUP0_AOI21X11_A_F_Z_R_10 0.1
`define C12T32_LLUP0_AOI21X11_B_R_Z_F_10 0.1
`define C12T32_LLUP0_AOI21X11_B_F_Z_R_10 0.1
`define C12T32_LLUP0_AOI21X11_C_R_Z_F_00 0.1
`define C12T32_LLUP0_AOI21X11_C_F_Z_R_00 0.1
`define C12T32_LLUP0_AOI21X11_C_R_Z_F_10 0.1
`define C12T32_LLUP0_AOI21X11_C_F_Z_R_10 0.1
`define C12T32_LLUP0_AOI21X11_C_R_Z_F_01 0.1
`define C12T32_LLUP0_AOI21X11_C_F_Z_R_01 0.1

module C12T32_LLUP0_AOI21X11 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL2, A, B) ;
	or    U2 (INTERNAL1, INTERNAL2, C) ;
	not   #1 U3 (Z, INTERNAL1) ;



	specify

		if (B && !C) (A -=> Z) = (`C12T32_LLUP0_AOI21X11_A_F_Z_R_10,`C12T32_LLUP0_AOI21X11_A_R_Z_F_10);
		if (A && !C) (B -=> Z) = (`C12T32_LLUP0_AOI21X11_B_F_Z_R_10,`C12T32_LLUP0_AOI21X11_B_R_Z_F_10);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_AOI21X11_C_F_Z_R_00,`C12T32_LLUP0_AOI21X11_C_R_Z_F_00);
		if (A && !B) (C -=> Z) = (`C12T32_LLUP0_AOI21X11_C_F_Z_R_10,`C12T32_LLUP0_AOI21X11_C_R_Z_F_10);
		if (!A && B) (C -=> Z) = (`C12T32_LLUP0_AOI21X11_C_F_Z_R_01,`C12T32_LLUP0_AOI21X11_C_R_Z_F_01);


	endspecify

endmodule // C12T32_LLUP0_AOI21X11


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_BFX134_A_R_Z_R 0.1
`define C12T32_LLUP0_BFX134_A_F_Z_F 0.1

module C12T32_LLUP0_BFX134 (Z, A);

	output Z;
	input A;

	buf   #1 U1 (Z, A) ;



	specify

		(A +=> Z) = (`C12T32_LLUP0_BFX134_A_R_Z_R,`C12T32_LLUP0_BFX134_A_F_Z_F);


	endspecify

endmodule // C12T32_LLUP0_BFX134


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_BFX16_A_R_Z_R 0.1
`define C12T32_LLUP0_BFX16_A_F_Z_F 0.1

module C12T32_LLUP0_BFX16 (Z, A);

	output Z;
	input A;

	buf   #1 U1 (Z, A) ;



	specify

		(A +=> Z) = (`C12T32_LLUP0_BFX16_A_R_Z_R,`C12T32_LLUP0_BFX16_A_F_Z_F);


	endspecify

endmodule // C12T32_LLUP0_BFX16


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_BFX33_A_R_Z_R 0.1
`define C12T32_LLUP0_BFX33_A_F_Z_F 0.1

module C12T32_LLUP0_BFX33 (Z, A);

	output Z;
	input A;

	buf   #1 U1 (Z, A) ;



	specify

		(A +=> Z) = (`C12T32_LLUP0_BFX33_A_R_Z_R,`C12T32_LLUP0_BFX33_A_F_Z_F);


	endspecify

endmodule // C12T32_LLUP0_BFX33


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_BFX4_A_R_Z_R 0.1
`define C12T32_LLUP0_BFX4_A_F_Z_F 0.1

module C12T32_LLUP0_BFX4 (Z, A);

	output Z;
	input A;

	buf   #1 U1 (Z, A) ;



	specify

		(A +=> Z) = (`C12T32_LLUP0_BFX4_A_R_Z_R,`C12T32_LLUP0_BFX4_A_F_Z_F);


	endspecify

endmodule // C12T32_LLUP0_BFX4


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_BFX67_A_R_Z_R 0.1
`define C12T32_LLUP0_BFX67_A_F_Z_F 0.1

module C12T32_LLUP0_BFX67 (Z, A);

	output Z;
	input A;

	buf   #1 U1 (Z, A) ;



	specify

		(A +=> Z) = (`C12T32_LLUP0_BFX67_A_R_Z_R,`C12T32_LLUP0_BFX67_A_F_Z_F);


	endspecify

endmodule // C12T32_LLUP0_BFX67


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_BFX8_A_R_Z_R 0.1
`define C12T32_LLUP0_BFX8_A_F_Z_F 0.1

module C12T32_LLUP0_BFX8 (Z, A);

	output Z;
	input A;

	buf   #1 U1 (Z, A) ;



	specify

		(A +=> Z) = (`C12T32_LLUP0_BFX8_A_R_Z_R,`C12T32_LLUP0_BFX8_A_F_Z_F);


	endspecify

endmodule // C12T32_LLUP0_BFX8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_CBI4I6X11_A_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X11_A_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X11_B_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X11_B_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X11_C_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X11_C_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X11_C_R_Z_F_110 0.1
`define C12T32_LLUP0_CBI4I6X11_C_F_Z_R_110 0.1
`define C12T32_LLUP0_CBI4I6X11_C_R_Z_F_100 0.1
`define C12T32_LLUP0_CBI4I6X11_C_F_Z_R_100 0.1
`define C12T32_LLUP0_CBI4I6X11_D_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X11_D_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X11_D_R_Z_F_001 0.1
`define C12T32_LLUP0_CBI4I6X11_D_F_Z_R_001 0.1
`define C12T32_LLUP0_CBI4I6X11_D_R_Z_F_000 0.1
`define C12T32_LLUP0_CBI4I6X11_D_F_Z_R_000 0.1
`define C12T32_LLUP0_CBI4I6X11_D_R_Z_F_110 0.1
`define C12T32_LLUP0_CBI4I6X11_D_F_Z_R_110 0.1
`define C12T32_LLUP0_CBI4I6X11_D_R_Z_F_100 0.1
`define C12T32_LLUP0_CBI4I6X11_D_F_Z_R_100 0.1

module C12T32_LLUP0_CBI4I6X11 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	or    U1 (INTERNAL3, A, B) ;
	and    U2 (INTERNAL2, INTERNAL3, C) ;
	or    U3 (INTERNAL1, INTERNAL2, D) ;
	not   #1 U4 (Z, INTERNAL1) ;



	specify

		if (!B && C && !D) (A -=> Z) = (`C12T32_LLUP0_CBI4I6X11_A_F_Z_R_010,`C12T32_LLUP0_CBI4I6X11_A_R_Z_F_010);
		if (!A && C && !D) (B -=> Z) = (`C12T32_LLUP0_CBI4I6X11_B_F_Z_R_010,`C12T32_LLUP0_CBI4I6X11_B_R_Z_F_010);
		if (!A && B && !D) (C -=> Z) = (`C12T32_LLUP0_CBI4I6X11_C_F_Z_R_010,`C12T32_LLUP0_CBI4I6X11_C_R_Z_F_010);
		if (A && B && !D) (C -=> Z) = (`C12T32_LLUP0_CBI4I6X11_C_F_Z_R_110,`C12T32_LLUP0_CBI4I6X11_C_R_Z_F_110);
		if (A && !B && !D) (C -=> Z) = (`C12T32_LLUP0_CBI4I6X11_C_F_Z_R_100,`C12T32_LLUP0_CBI4I6X11_C_R_Z_F_100);
		if (!A && B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X11_D_F_Z_R_010,`C12T32_LLUP0_CBI4I6X11_D_R_Z_F_010);
		if (!A && !B && C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X11_D_F_Z_R_001,`C12T32_LLUP0_CBI4I6X11_D_R_Z_F_001);
		if (!A && !B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X11_D_F_Z_R_000,`C12T32_LLUP0_CBI4I6X11_D_R_Z_F_000);
		if (A && B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X11_D_F_Z_R_110,`C12T32_LLUP0_CBI4I6X11_D_R_Z_F_110);
		if (A && !B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X11_D_F_Z_R_100,`C12T32_LLUP0_CBI4I6X11_D_R_Z_F_100);


	endspecify

endmodule // C12T32_LLUP0_CBI4I6X11


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_CBI4I6X5_A_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X5_A_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X5_B_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X5_B_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X5_C_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X5_C_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X5_C_R_Z_F_110 0.1
`define C12T32_LLUP0_CBI4I6X5_C_F_Z_R_110 0.1
`define C12T32_LLUP0_CBI4I6X5_C_R_Z_F_100 0.1
`define C12T32_LLUP0_CBI4I6X5_C_F_Z_R_100 0.1
`define C12T32_LLUP0_CBI4I6X5_D_R_Z_F_010 0.1
`define C12T32_LLUP0_CBI4I6X5_D_F_Z_R_010 0.1
`define C12T32_LLUP0_CBI4I6X5_D_R_Z_F_001 0.1
`define C12T32_LLUP0_CBI4I6X5_D_F_Z_R_001 0.1
`define C12T32_LLUP0_CBI4I6X5_D_R_Z_F_000 0.1
`define C12T32_LLUP0_CBI4I6X5_D_F_Z_R_000 0.1
`define C12T32_LLUP0_CBI4I6X5_D_R_Z_F_110 0.1
`define C12T32_LLUP0_CBI4I6X5_D_F_Z_R_110 0.1
`define C12T32_LLUP0_CBI4I6X5_D_R_Z_F_100 0.1
`define C12T32_LLUP0_CBI4I6X5_D_F_Z_R_100 0.1

module C12T32_LLUP0_CBI4I6X5 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	or    U1 (INTERNAL3, A, B) ;
	and    U2 (INTERNAL2, INTERNAL3, C) ;
	or    U3 (INTERNAL1, INTERNAL2, D) ;
	not   #1 U4 (Z, INTERNAL1) ;



	specify

		if (!B && C && !D) (A -=> Z) = (`C12T32_LLUP0_CBI4I6X5_A_F_Z_R_010,`C12T32_LLUP0_CBI4I6X5_A_R_Z_F_010);
		if (!A && C && !D) (B -=> Z) = (`C12T32_LLUP0_CBI4I6X5_B_F_Z_R_010,`C12T32_LLUP0_CBI4I6X5_B_R_Z_F_010);
		if (!A && B && !D) (C -=> Z) = (`C12T32_LLUP0_CBI4I6X5_C_F_Z_R_010,`C12T32_LLUP0_CBI4I6X5_C_R_Z_F_010);
		if (A && B && !D) (C -=> Z) = (`C12T32_LLUP0_CBI4I6X5_C_F_Z_R_110,`C12T32_LLUP0_CBI4I6X5_C_R_Z_F_110);
		if (A && !B && !D) (C -=> Z) = (`C12T32_LLUP0_CBI4I6X5_C_F_Z_R_100,`C12T32_LLUP0_CBI4I6X5_C_R_Z_F_100);
		if (!A && B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X5_D_F_Z_R_010,`C12T32_LLUP0_CBI4I6X5_D_R_Z_F_010);
		if (!A && !B && C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X5_D_F_Z_R_001,`C12T32_LLUP0_CBI4I6X5_D_R_Z_F_001);
		if (!A && !B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X5_D_F_Z_R_000,`C12T32_LLUP0_CBI4I6X5_D_R_Z_F_000);
		if (A && B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X5_D_F_Z_R_110,`C12T32_LLUP0_CBI4I6X5_D_R_Z_F_110);
		if (A && !B && !C) (D -=> Z) = (`C12T32_LLUP0_CBI4I6X5_D_F_Z_R_100,`C12T32_LLUP0_CBI4I6X5_D_R_Z_F_100);


	endspecify

endmodule // C12T32_LLUP0_CBI4I6X5


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_FA1X6_A0_R_CO_R_10 0.1
`define C12T32_LLUP0_FA1X6_A0_F_CO_F_10 0.1
`define C12T32_LLUP0_FA1X6_A0_R_CO_R_01 0.1
`define C12T32_LLUP0_FA1X6_A0_F_CO_F_01 0.1
`define C12T32_LLUP0_FA1X6_A0_R_S0_F_10 0.1
`define C12T32_LLUP0_FA1X6_A0_F_S0_R_10 0.1
`define C12T32_LLUP0_FA1X6_A0_R_S0_F_01 0.1
`define C12T32_LLUP0_FA1X6_A0_F_S0_R_01 0.1
`define C12T32_LLUP0_FA1X6_A0_R_S0_R_00 0.1
`define C12T32_LLUP0_FA1X6_A0_F_S0_F_00 0.1
`define C12T32_LLUP0_FA1X6_A0_R_S0_R_11 0.1
`define C12T32_LLUP0_FA1X6_A0_F_S0_F_11 0.1
`define C12T32_LLUP0_FA1X6_B0_R_CO_R_10 0.1
`define C12T32_LLUP0_FA1X6_B0_F_CO_F_10 0.1
`define C12T32_LLUP0_FA1X6_B0_R_CO_R_01 0.1
`define C12T32_LLUP0_FA1X6_B0_F_CO_F_01 0.1
`define C12T32_LLUP0_FA1X6_B0_R_S0_F_10 0.1
`define C12T32_LLUP0_FA1X6_B0_F_S0_R_10 0.1
`define C12T32_LLUP0_FA1X6_B0_R_S0_F_01 0.1
`define C12T32_LLUP0_FA1X6_B0_F_S0_R_01 0.1
`define C12T32_LLUP0_FA1X6_B0_R_S0_R_00 0.1
`define C12T32_LLUP0_FA1X6_B0_F_S0_F_00 0.1
`define C12T32_LLUP0_FA1X6_B0_R_S0_R_11 0.1
`define C12T32_LLUP0_FA1X6_B0_F_S0_F_11 0.1
`define C12T32_LLUP0_FA1X6_CI_R_CO_R_10 0.1
`define C12T32_LLUP0_FA1X6_CI_F_CO_F_10 0.1
`define C12T32_LLUP0_FA1X6_CI_R_CO_R_01 0.1
`define C12T32_LLUP0_FA1X6_CI_F_CO_F_01 0.1
`define C12T32_LLUP0_FA1X6_CI_R_S0_F_10 0.1
`define C12T32_LLUP0_FA1X6_CI_F_S0_R_10 0.1
`define C12T32_LLUP0_FA1X6_CI_R_S0_F_01 0.1
`define C12T32_LLUP0_FA1X6_CI_F_S0_R_01 0.1
`define C12T32_LLUP0_FA1X6_CI_R_S0_R_00 0.1
`define C12T32_LLUP0_FA1X6_CI_F_S0_F_00 0.1
`define C12T32_LLUP0_FA1X6_CI_R_S0_R_11 0.1
`define C12T32_LLUP0_FA1X6_CI_F_S0_F_11 0.1

module C12T32_LLUP0_FA1X6 (S0, CO, A0, B0, CI);

	output S0;
	output CO;
	input A0;
	input B0;
	input CI;

	xor   #1 U1 (S0, A0, B0, CI) ;
	or    U2 (INTERNAL2, A0, B0) ;
	and    U3 (INTERNAL1, INTERNAL2, CI) ;
	and    U4 (INTERNAL3, A0, B0) ;
	or   #1 U5 (CO, INTERNAL1, INTERNAL3) ;



	specify

		if (B0 && !CI) (A0 +=> CO) = (`C12T32_LLUP0_FA1X6_A0_R_CO_R_10,`C12T32_LLUP0_FA1X6_A0_F_CO_F_10);
		if (!B0 && CI) (A0 +=> CO) = (`C12T32_LLUP0_FA1X6_A0_R_CO_R_01,`C12T32_LLUP0_FA1X6_A0_F_CO_F_01);
		if (B0 && !CI) (A0 -=> S0) = (`C12T32_LLUP0_FA1X6_A0_F_S0_R_10,`C12T32_LLUP0_FA1X6_A0_R_S0_F_10);
		if (!B0 && CI) (A0 -=> S0) = (`C12T32_LLUP0_FA1X6_A0_F_S0_R_01,`C12T32_LLUP0_FA1X6_A0_R_S0_F_01);
		if (!B0 && !CI) (A0 +=> S0) = (`C12T32_LLUP0_FA1X6_A0_R_S0_R_00,`C12T32_LLUP0_FA1X6_A0_F_S0_F_00);
		if (B0 && CI) (A0 +=> S0) = (`C12T32_LLUP0_FA1X6_A0_R_S0_R_11,`C12T32_LLUP0_FA1X6_A0_F_S0_F_11);
		if (A0 && !CI) (B0 +=> CO) = (`C12T32_LLUP0_FA1X6_B0_R_CO_R_10,`C12T32_LLUP0_FA1X6_B0_F_CO_F_10);
		if (!A0 && CI) (B0 +=> CO) = (`C12T32_LLUP0_FA1X6_B0_R_CO_R_01,`C12T32_LLUP0_FA1X6_B0_F_CO_F_01);
		if (A0 && !CI) (B0 -=> S0) = (`C12T32_LLUP0_FA1X6_B0_F_S0_R_10,`C12T32_LLUP0_FA1X6_B0_R_S0_F_10);
		if (!A0 && CI) (B0 -=> S0) = (`C12T32_LLUP0_FA1X6_B0_F_S0_R_01,`C12T32_LLUP0_FA1X6_B0_R_S0_F_01);
		if (!A0 && !CI) (B0 +=> S0) = (`C12T32_LLUP0_FA1X6_B0_R_S0_R_00,`C12T32_LLUP0_FA1X6_B0_F_S0_F_00);
		if (A0 && CI) (B0 +=> S0) = (`C12T32_LLUP0_FA1X6_B0_R_S0_R_11,`C12T32_LLUP0_FA1X6_B0_F_S0_F_11);
		if (A0 && !B0) (CI +=> CO) = (`C12T32_LLUP0_FA1X6_CI_R_CO_R_10,`C12T32_LLUP0_FA1X6_CI_F_CO_F_10);
		if (!A0 && B0) (CI +=> CO) = (`C12T32_LLUP0_FA1X6_CI_R_CO_R_01,`C12T32_LLUP0_FA1X6_CI_F_CO_F_01);
		if (A0 && !B0) (CI -=> S0) = (`C12T32_LLUP0_FA1X6_CI_F_S0_R_10,`C12T32_LLUP0_FA1X6_CI_R_S0_F_10);
		if (!A0 && B0) (CI -=> S0) = (`C12T32_LLUP0_FA1X6_CI_F_S0_R_01,`C12T32_LLUP0_FA1X6_CI_R_S0_F_01);
		if (!A0 && !B0) (CI +=> S0) = (`C12T32_LLUP0_FA1X6_CI_R_S0_R_00,`C12T32_LLUP0_FA1X6_CI_F_S0_F_00);
		if (A0 && B0) (CI +=> S0) = (`C12T32_LLUP0_FA1X6_CI_R_S0_R_11,`C12T32_LLUP0_FA1X6_CI_F_S0_F_11);


	endspecify

endmodule // C12T32_LLUP0_FA1X6


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_FA1X8_A0_R_CO_R_10 0.1
`define C12T32_LLUP0_FA1X8_A0_F_CO_F_10 0.1
`define C12T32_LLUP0_FA1X8_A0_R_CO_R_01 0.1
`define C12T32_LLUP0_FA1X8_A0_F_CO_F_01 0.1
`define C12T32_LLUP0_FA1X8_A0_R_S0_F_10 0.1
`define C12T32_LLUP0_FA1X8_A0_F_S0_R_10 0.1
`define C12T32_LLUP0_FA1X8_A0_R_S0_F_01 0.1
`define C12T32_LLUP0_FA1X8_A0_F_S0_R_01 0.1
`define C12T32_LLUP0_FA1X8_A0_R_S0_R_00 0.1
`define C12T32_LLUP0_FA1X8_A0_F_S0_F_00 0.1
`define C12T32_LLUP0_FA1X8_A0_R_S0_R_11 0.1
`define C12T32_LLUP0_FA1X8_A0_F_S0_F_11 0.1
`define C12T32_LLUP0_FA1X8_B0_R_CO_R_10 0.1
`define C12T32_LLUP0_FA1X8_B0_F_CO_F_10 0.1
`define C12T32_LLUP0_FA1X8_B0_R_CO_R_01 0.1
`define C12T32_LLUP0_FA1X8_B0_F_CO_F_01 0.1
`define C12T32_LLUP0_FA1X8_B0_R_S0_F_10 0.1
`define C12T32_LLUP0_FA1X8_B0_F_S0_R_10 0.1
`define C12T32_LLUP0_FA1X8_B0_R_S0_F_01 0.1
`define C12T32_LLUP0_FA1X8_B0_F_S0_R_01 0.1
`define C12T32_LLUP0_FA1X8_B0_R_S0_R_00 0.1
`define C12T32_LLUP0_FA1X8_B0_F_S0_F_00 0.1
`define C12T32_LLUP0_FA1X8_B0_R_S0_R_11 0.1
`define C12T32_LLUP0_FA1X8_B0_F_S0_F_11 0.1
`define C12T32_LLUP0_FA1X8_CI_R_CO_R_10 0.1
`define C12T32_LLUP0_FA1X8_CI_F_CO_F_10 0.1
`define C12T32_LLUP0_FA1X8_CI_R_CO_R_01 0.1
`define C12T32_LLUP0_FA1X8_CI_F_CO_F_01 0.1
`define C12T32_LLUP0_FA1X8_CI_R_S0_F_10 0.1
`define C12T32_LLUP0_FA1X8_CI_F_S0_R_10 0.1
`define C12T32_LLUP0_FA1X8_CI_R_S0_F_01 0.1
`define C12T32_LLUP0_FA1X8_CI_F_S0_R_01 0.1
`define C12T32_LLUP0_FA1X8_CI_R_S0_R_00 0.1
`define C12T32_LLUP0_FA1X8_CI_F_S0_F_00 0.1
`define C12T32_LLUP0_FA1X8_CI_R_S0_R_11 0.1
`define C12T32_LLUP0_FA1X8_CI_F_S0_F_11 0.1

module C12T32_LLUP0_FA1X8 (S0, CO, A0, B0, CI);

	output S0;
	output CO;
	input A0;
	input B0;
	input CI;

	xor   #1 U1 (S0, A0, B0, CI) ;
	or    U2 (INTERNAL2, A0, B0) ;
	and    U3 (INTERNAL1, INTERNAL2, CI) ;
	and    U4 (INTERNAL3, A0, B0) ;
	or   #1 U5 (CO, INTERNAL1, INTERNAL3) ;



	specify

		if (B0 && !CI) (A0 +=> CO) = (`C12T32_LLUP0_FA1X8_A0_R_CO_R_10,`C12T32_LLUP0_FA1X8_A0_F_CO_F_10);
		if (!B0 && CI) (A0 +=> CO) = (`C12T32_LLUP0_FA1X8_A0_R_CO_R_01,`C12T32_LLUP0_FA1X8_A0_F_CO_F_01);
		if (B0 && !CI) (A0 -=> S0) = (`C12T32_LLUP0_FA1X8_A0_F_S0_R_10,`C12T32_LLUP0_FA1X8_A0_R_S0_F_10);
		if (!B0 && CI) (A0 -=> S0) = (`C12T32_LLUP0_FA1X8_A0_F_S0_R_01,`C12T32_LLUP0_FA1X8_A0_R_S0_F_01);
		if (!B0 && !CI) (A0 +=> S0) = (`C12T32_LLUP0_FA1X8_A0_R_S0_R_00,`C12T32_LLUP0_FA1X8_A0_F_S0_F_00);
		if (B0 && CI) (A0 +=> S0) = (`C12T32_LLUP0_FA1X8_A0_R_S0_R_11,`C12T32_LLUP0_FA1X8_A0_F_S0_F_11);
		if (A0 && !CI) (B0 +=> CO) = (`C12T32_LLUP0_FA1X8_B0_R_CO_R_10,`C12T32_LLUP0_FA1X8_B0_F_CO_F_10);
		if (!A0 && CI) (B0 +=> CO) = (`C12T32_LLUP0_FA1X8_B0_R_CO_R_01,`C12T32_LLUP0_FA1X8_B0_F_CO_F_01);
		if (A0 && !CI) (B0 -=> S0) = (`C12T32_LLUP0_FA1X8_B0_F_S0_R_10,`C12T32_LLUP0_FA1X8_B0_R_S0_F_10);
		if (!A0 && CI) (B0 -=> S0) = (`C12T32_LLUP0_FA1X8_B0_F_S0_R_01,`C12T32_LLUP0_FA1X8_B0_R_S0_F_01);
		if (!A0 && !CI) (B0 +=> S0) = (`C12T32_LLUP0_FA1X8_B0_R_S0_R_00,`C12T32_LLUP0_FA1X8_B0_F_S0_F_00);
		if (A0 && CI) (B0 +=> S0) = (`C12T32_LLUP0_FA1X8_B0_R_S0_R_11,`C12T32_LLUP0_FA1X8_B0_F_S0_F_11);
		if (A0 && !B0) (CI +=> CO) = (`C12T32_LLUP0_FA1X8_CI_R_CO_R_10,`C12T32_LLUP0_FA1X8_CI_F_CO_F_10);
		if (!A0 && B0) (CI +=> CO) = (`C12T32_LLUP0_FA1X8_CI_R_CO_R_01,`C12T32_LLUP0_FA1X8_CI_F_CO_F_01);
		if (A0 && !B0) (CI -=> S0) = (`C12T32_LLUP0_FA1X8_CI_F_S0_R_10,`C12T32_LLUP0_FA1X8_CI_R_S0_F_10);
		if (!A0 && B0) (CI -=> S0) = (`C12T32_LLUP0_FA1X8_CI_F_S0_R_01,`C12T32_LLUP0_FA1X8_CI_R_S0_F_01);
		if (!A0 && !B0) (CI +=> S0) = (`C12T32_LLUP0_FA1X8_CI_R_S0_R_00,`C12T32_LLUP0_FA1X8_CI_F_S0_F_00);
		if (A0 && B0) (CI +=> S0) = (`C12T32_LLUP0_FA1X8_CI_R_S0_R_11,`C12T32_LLUP0_FA1X8_CI_F_S0_F_11);


	endspecify

endmodule // C12T32_LLUP0_FA1X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_IVX134_A_R_Z_F 0.1
`define C12T32_LLUP0_IVX134_A_F_Z_R 0.1

module C12T32_LLUP0_IVX134 (Z, A);

	output Z;
	input A;

	not   #1 U1 (Z, A) ;



	specify

		(A -=> Z) = (`C12T32_LLUP0_IVX134_A_F_Z_R,`C12T32_LLUP0_IVX134_A_R_Z_F);


	endspecify

endmodule // C12T32_LLUP0_IVX134


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_IVX17_A_R_Z_F 0.1
`define C12T32_LLUP0_IVX17_A_F_Z_R 0.1

module C12T32_LLUP0_IVX17 (Z, A);

	output Z;
	input A;

	not   #1 U1 (Z, A) ;



	specify

		(A -=> Z) = (`C12T32_LLUP0_IVX17_A_F_Z_R,`C12T32_LLUP0_IVX17_A_R_Z_F);


	endspecify

endmodule // C12T32_LLUP0_IVX17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_IVX33_A_R_Z_F 0.1
`define C12T32_LLUP0_IVX33_A_F_Z_R 0.1

module C12T32_LLUP0_IVX33 (Z, A);

	output Z;
	input A;

	not   #1 U1 (Z, A) ;



	specify

		(A -=> Z) = (`C12T32_LLUP0_IVX33_A_F_Z_R,`C12T32_LLUP0_IVX33_A_R_Z_F);


	endspecify

endmodule // C12T32_LLUP0_IVX33


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_IVX4_A_R_Z_F 0.1
`define C12T32_LLUP0_IVX4_A_F_Z_R 0.1

module C12T32_LLUP0_IVX4 (Z, A);

	output Z;
	input A;

	not   #1 U1 (Z, A) ;



	specify

		(A -=> Z) = (`C12T32_LLUP0_IVX4_A_F_Z_R,`C12T32_LLUP0_IVX4_A_R_Z_F);


	endspecify

endmodule // C12T32_LLUP0_IVX4


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_IVX67_A_R_Z_F 0.1
`define C12T32_LLUP0_IVX67_A_F_Z_R 0.1

module C12T32_LLUP0_IVX67 (Z, A);

	output Z;
	input A;

	not   #1 U1 (Z, A) ;



	specify

		(A -=> Z) = (`C12T32_LLUP0_IVX67_A_F_Z_R,`C12T32_LLUP0_IVX67_A_R_Z_F);


	endspecify

endmodule // C12T32_LLUP0_IVX67


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_IVX8_A_R_Z_F 0.1
`define C12T32_LLUP0_IVX8_A_F_Z_R 0.1

module C12T32_LLUP0_IVX8 (Z, A);

	output Z;
	input A;

	not   #1 U1 (Z, A) ;



	specify

		(A -=> Z) = (`C12T32_LLUP0_IVX8_A_F_Z_R,`C12T32_LLUP0_IVX8_A_R_Z_F);


	endspecify

endmodule // C12T32_LLUP0_IVX8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUX21X17_D0_R_Z_R_00 0.1
`define C12T32_LLUP0_MUX21X17_D0_F_Z_F_00 0.1
`define C12T32_LLUP0_MUX21X17_D0_R_Z_R_10 0.1
`define C12T32_LLUP0_MUX21X17_D0_F_Z_F_10 0.1
`define C12T32_LLUP0_MUX21X17_D1_R_Z_R_01 0.1
`define C12T32_LLUP0_MUX21X17_D1_F_Z_F_01 0.1
`define C12T32_LLUP0_MUX21X17_D1_R_Z_R_11 0.1
`define C12T32_LLUP0_MUX21X17_D1_F_Z_F_11 0.1
`define C12T32_LLUP0_MUX21X17_S0_R_Z_F_10 0.1
`define C12T32_LLUP0_MUX21X17_S0_F_Z_R_10 0.1
`define C12T32_LLUP0_MUX21X17_S0_R_Z_R_01 0.1
`define C12T32_LLUP0_MUX21X17_S0_F_Z_F_01 0.1

module C12T32_LLUP0_MUX21X17 (Z, D0, D1, S0);

	output Z;
	input D0;
	input D1;
	input S0;

	U_MUX2  #1 U1 (Z, D0, D1, S0) ;



	specify

		if (!D1 && !S0) (D0 +=> Z) = (`C12T32_LLUP0_MUX21X17_D0_R_Z_R_00,`C12T32_LLUP0_MUX21X17_D0_F_Z_F_00);
		if (D1 && !S0) (D0 +=> Z) = (`C12T32_LLUP0_MUX21X17_D0_R_Z_R_10,`C12T32_LLUP0_MUX21X17_D0_F_Z_F_10);
		if (!D0 && S0) (D1 +=> Z) = (`C12T32_LLUP0_MUX21X17_D1_R_Z_R_01,`C12T32_LLUP0_MUX21X17_D1_F_Z_F_01);
		if (D0 && S0) (D1 +=> Z) = (`C12T32_LLUP0_MUX21X17_D1_R_Z_R_11,`C12T32_LLUP0_MUX21X17_D1_F_Z_F_11);
		if (D0 && !D1) (S0 -=> Z) = (`C12T32_LLUP0_MUX21X17_S0_F_Z_R_10,`C12T32_LLUP0_MUX21X17_S0_R_Z_F_10);
		if (!D0 && D1) (S0 +=> Z) = (`C12T32_LLUP0_MUX21X17_S0_R_Z_R_01,`C12T32_LLUP0_MUX21X17_S0_F_Z_F_01);


	endspecify

endmodule // C12T32_LLUP0_MUX21X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUX21X8_D0_R_Z_R_00 0.1
`define C12T32_LLUP0_MUX21X8_D0_F_Z_F_00 0.1
`define C12T32_LLUP0_MUX21X8_D0_R_Z_R_10 0.1
`define C12T32_LLUP0_MUX21X8_D0_F_Z_F_10 0.1
`define C12T32_LLUP0_MUX21X8_D1_R_Z_R_01 0.1
`define C12T32_LLUP0_MUX21X8_D1_F_Z_F_01 0.1
`define C12T32_LLUP0_MUX21X8_D1_R_Z_R_11 0.1
`define C12T32_LLUP0_MUX21X8_D1_F_Z_F_11 0.1
`define C12T32_LLUP0_MUX21X8_S0_R_Z_F_10 0.1
`define C12T32_LLUP0_MUX21X8_S0_F_Z_R_10 0.1
`define C12T32_LLUP0_MUX21X8_S0_R_Z_R_01 0.1
`define C12T32_LLUP0_MUX21X8_S0_F_Z_F_01 0.1

module C12T32_LLUP0_MUX21X8 (Z, D0, D1, S0);

	output Z;
	input D0;
	input D1;
	input S0;

	U_MUX2  #1 U1 (Z, D0, D1, S0) ;



	specify

		if (!D1 && !S0) (D0 +=> Z) = (`C12T32_LLUP0_MUX21X8_D0_R_Z_R_00,`C12T32_LLUP0_MUX21X8_D0_F_Z_F_00);
		if (D1 && !S0) (D0 +=> Z) = (`C12T32_LLUP0_MUX21X8_D0_R_Z_R_10,`C12T32_LLUP0_MUX21X8_D0_F_Z_F_10);
		if (!D0 && S0) (D1 +=> Z) = (`C12T32_LLUP0_MUX21X8_D1_R_Z_R_01,`C12T32_LLUP0_MUX21X8_D1_F_Z_F_01);
		if (D0 && S0) (D1 +=> Z) = (`C12T32_LLUP0_MUX21X8_D1_R_Z_R_11,`C12T32_LLUP0_MUX21X8_D1_F_Z_F_11);
		if (D0 && !D1) (S0 -=> Z) = (`C12T32_LLUP0_MUX21X8_S0_F_Z_R_10,`C12T32_LLUP0_MUX21X8_S0_R_Z_F_10);
		if (!D0 && D1) (S0 +=> Z) = (`C12T32_LLUP0_MUX21X8_S0_R_Z_R_01,`C12T32_LLUP0_MUX21X8_S0_F_Z_F_01);


	endspecify

endmodule // C12T32_LLUP0_MUX21X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_00000 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_00000 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_10100 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_10100 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_11000 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_11000 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_11100 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_11100 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_10000 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_10000 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_00100 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_00100 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_01000 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_01000 0.1
`define C12T32_LLUP0_MUX41X31_D0_R_Z_R_01100 0.1
`define C12T32_LLUP0_MUX41X31_D0_F_Z_F_01100 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_00010 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_00010 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_10110 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_10110 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_11010 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_11010 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_11110 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_11110 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_10010 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_10010 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_00110 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_00110 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_01010 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_01010 0.1
`define C12T32_LLUP0_MUX41X31_D1_R_Z_R_01110 0.1
`define C12T32_LLUP0_MUX41X31_D1_F_Z_F_01110 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_00001 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_00001 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_10101 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_10101 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_11001 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_11001 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_11101 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_11101 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_10001 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_10001 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_00101 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_00101 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_01001 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_01001 0.1
`define C12T32_LLUP0_MUX41X31_D2_R_Z_R_01101 0.1
`define C12T32_LLUP0_MUX41X31_D2_F_Z_F_01101 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_00011 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_00011 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_10111 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_10111 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_11011 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_11011 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_11111 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_11111 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_10011 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_10011 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_00111 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_00111 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_01011 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_01011 0.1
`define C12T32_LLUP0_MUX41X31_D3_R_Z_R_01111 0.1
`define C12T32_LLUP0_MUX41X31_D3_F_Z_F_01111 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_00101 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_00101 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_10101 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_10101 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_10110 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_10110 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_11101 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_11101 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_10100 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_10100 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_01101 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_01101 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_10000 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_10000 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_F_10010 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_R_10010 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_00011 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_00011 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_01110 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_01110 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_10011 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_10011 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_11011 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_11011 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_01100 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_01100 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_01000 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_01000 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_01010 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_01010 0.1
`define C12T32_LLUP0_MUX41X31_S0_R_Z_R_01011 0.1
`define C12T32_LLUP0_MUX41X31_S0_F_Z_F_01011 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_01001 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_01001 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_11001 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_11001 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_11010 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_11010 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_11101 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_11101 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_11000 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_11000 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_01101 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_01101 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_10000 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_10000 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_F_10010 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_R_10010 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_00011 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_00011 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_01110 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_01110 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_10011 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_10011 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_10111 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_10111 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_01100 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_01100 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_00100 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_00100 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_00110 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_00110 0.1
`define C12T32_LLUP0_MUX41X31_S1_R_Z_R_00111 0.1
`define C12T32_LLUP0_MUX41X31_S1_F_Z_F_00111 0.1

module C12T32_LLUP0_MUX41X31 (Z, D0, D1, D2, D3, S0, S1);

	output Z;
	input D0;
	input D1;
	input D2;
	input D3;
	input S0;
	input S1;

	U_MUX2   U1 (INTERNAL1, D0, D1, S0) ;
	U_MUX2   U2 (INTERNAL2, D2, D3, S0) ;
	U_MUX2  #1 U3 (Z, INTERNAL1, INTERNAL2, S1) ;



	specify

		if (!D1 && !D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_00000,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_00000);
		if (D1 && !D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_10100,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_10100);
		if (D1 && D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_11000,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_11000);
		if (D1 && D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_11100,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_11100);
		if (D1 && !D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_10000,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_10000);
		if (!D1 && !D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_00100,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_00100);
		if (!D1 && D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_01000,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_01000);
		if (!D1 && D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X31_D0_R_Z_R_01100,`C12T32_LLUP0_MUX41X31_D0_F_Z_F_01100);
		if (!D0 && !D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_00010,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_00010);
		if (D0 && !D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_10110,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_10110);
		if (D0 && D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_11010,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_11010);
		if (D0 && D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_11110,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_11110);
		if (D0 && !D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_10010,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_10010);
		if (!D0 && !D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_00110,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_00110);
		if (!D0 && D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_01010,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_01010);
		if (!D0 && D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X31_D1_R_Z_R_01110,`C12T32_LLUP0_MUX41X31_D1_F_Z_F_01110);
		if (!D0 && !D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_00001,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_00001);
		if (D0 && !D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_10101,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_10101);
		if (D0 && D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_11001,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_11001);
		if (D0 && D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_11101,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_11101);
		if (D0 && !D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_10001,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_10001);
		if (!D0 && !D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_00101,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_00101);
		if (!D0 && D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_01001,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_01001);
		if (!D0 && D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X31_D2_R_Z_R_01101,`C12T32_LLUP0_MUX41X31_D2_F_Z_F_01101);
		if (!D0 && !D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_00011,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_00011);
		if (D0 && !D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_10111,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_10111);
		if (D0 && D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_11011,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_11011);
		if (D0 && D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_11111,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_11111);
		if (D0 && !D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_10011,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_10011);
		if (!D0 && !D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_00111,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_00111);
		if (!D0 && D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_01011,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_01011);
		if (!D0 && D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X31_D3_R_Z_R_01111,`C12T32_LLUP0_MUX41X31_D3_F_Z_F_01111);
		if (!D0 && !D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_00101,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_00101);
		if (D0 && !D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_10101,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_10101);
		if (D0 && !D1 && D2 && D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_10110,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_10110);
		if (D0 && D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_11101,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_11101);
		if (D0 && !D1 && D2 && !D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_10100,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_10100);
		if (!D0 && D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_01101,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_01101);
		if (D0 && !D1 && !D2 && !D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_10000,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_10000);
		if (D0 && !D1 && !D2 && D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X31_S0_F_Z_R_10010,`C12T32_LLUP0_MUX41X31_S0_R_Z_F_10010);
		if (!D0 && !D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_00011,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_00011);
		if (!D0 && D1 && D2 && D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_01110,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_01110);
		if (D0 && !D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_10011,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_10011);
		if (D0 && D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_11011,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_11011);
		if (!D0 && D1 && D2 && !D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_01100,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_01100);
		if (!D0 && D1 && !D2 && !D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_01000,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_01000);
		if (!D0 && D1 && !D2 && D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_01010,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_01010);
		if (!D0 && D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X31_S0_R_Z_R_01011,`C12T32_LLUP0_MUX41X31_S0_F_Z_F_01011);
		if (!D0 && D1 && !D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_01001,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_01001);
		if (D0 && D1 && !D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_11001,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_11001);
		if (D0 && D1 && !D2 && D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_11010,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_11010);
		if (D0 && D1 && D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_11101,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_11101);
		if (D0 && D1 && !D2 && !D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_11000,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_11000);
		if (!D0 && D1 && D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_01101,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_01101);
		if (D0 && !D1 && !D2 && !D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_10000,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_10000);
		if (D0 && !D1 && !D2 && D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X31_S1_F_Z_R_10010,`C12T32_LLUP0_MUX41X31_S1_R_Z_F_10010);
		if (!D0 && !D1 && !D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_00011,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_00011);
		if (!D0 && D1 && D2 && D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_01110,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_01110);
		if (D0 && !D1 && !D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_10011,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_10011);
		if (D0 && !D1 && D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_10111,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_10111);
		if (!D0 && D1 && D2 && !D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_01100,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_01100);
		if (!D0 && !D1 && D2 && !D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_00100,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_00100);
		if (!D0 && !D1 && D2 && D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_00110,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_00110);
		if (!D0 && !D1 && D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X31_S1_R_Z_R_00111,`C12T32_LLUP0_MUX41X31_S1_F_Z_F_00111);


	endspecify

endmodule // C12T32_LLUP0_MUX41X31


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_00000 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_00000 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_10100 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_10100 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_11000 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_11000 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_11100 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_11100 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_10000 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_10000 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_00100 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_00100 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_01000 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_01000 0.1
`define C12T32_LLUP0_MUX41X8_D0_R_Z_R_01100 0.1
`define C12T32_LLUP0_MUX41X8_D0_F_Z_F_01100 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_00010 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_00010 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_10110 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_10110 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_11010 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_11010 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_11110 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_11110 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_10010 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_10010 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_00110 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_00110 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_01010 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_01010 0.1
`define C12T32_LLUP0_MUX41X8_D1_R_Z_R_01110 0.1
`define C12T32_LLUP0_MUX41X8_D1_F_Z_F_01110 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_00001 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_00001 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_10101 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_10101 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_11001 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_11001 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_11101 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_11101 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_10001 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_10001 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_00101 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_00101 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_01001 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_01001 0.1
`define C12T32_LLUP0_MUX41X8_D2_R_Z_R_01101 0.1
`define C12T32_LLUP0_MUX41X8_D2_F_Z_F_01101 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_00011 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_00011 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_10111 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_10111 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_11011 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_11011 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_11111 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_11111 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_10011 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_10011 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_00111 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_00111 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_01011 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_01011 0.1
`define C12T32_LLUP0_MUX41X8_D3_R_Z_R_01111 0.1
`define C12T32_LLUP0_MUX41X8_D3_F_Z_F_01111 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_00101 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_00101 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_10101 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_10101 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_10110 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_10110 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_11101 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_11101 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_10100 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_10100 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_01101 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_01101 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_10000 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_10000 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_F_10010 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_R_10010 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_00011 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_00011 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_01110 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_01110 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_10011 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_10011 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_11011 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_11011 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_01100 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_01100 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_01000 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_01000 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_01010 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_01010 0.1
`define C12T32_LLUP0_MUX41X8_S0_R_Z_R_01011 0.1
`define C12T32_LLUP0_MUX41X8_S0_F_Z_F_01011 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_01001 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_01001 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_11001 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_11001 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_11010 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_11010 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_11101 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_11101 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_11000 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_11000 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_01101 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_01101 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_10000 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_10000 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_F_10010 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_R_10010 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_00011 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_00011 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_01110 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_01110 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_10011 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_10011 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_10111 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_10111 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_01100 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_01100 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_00100 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_00100 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_00110 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_00110 0.1
`define C12T32_LLUP0_MUX41X8_S1_R_Z_R_00111 0.1
`define C12T32_LLUP0_MUX41X8_S1_F_Z_F_00111 0.1

module C12T32_LLUP0_MUX41X8 (Z, D0, D1, D2, D3, S0, S1);

	output Z;
	input D0;
	input D1;
	input D2;
	input D3;
	input S0;
	input S1;

	U_MUX2   U1 (INTERNAL1, D0, D1, S0) ;
	U_MUX2   U2 (INTERNAL2, D2, D3, S0) ;
	U_MUX2  #1 U3 (Z, INTERNAL1, INTERNAL2, S1) ;



	specify

		if (!D1 && !D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_00000,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_00000);
		if (D1 && !D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_10100,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_10100);
		if (D1 && D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_11000,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_11000);
		if (D1 && D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_11100,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_11100);
		if (D1 && !D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_10000,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_10000);
		if (!D1 && !D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_00100,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_00100);
		if (!D1 && D2 && !D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_01000,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_01000);
		if (!D1 && D2 && D3 && !S0 && !S1) (D0 +=> Z) = (`C12T32_LLUP0_MUX41X8_D0_R_Z_R_01100,`C12T32_LLUP0_MUX41X8_D0_F_Z_F_01100);
		if (!D0 && !D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_00010,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_00010);
		if (D0 && !D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_10110,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_10110);
		if (D0 && D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_11010,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_11010);
		if (D0 && D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_11110,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_11110);
		if (D0 && !D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_10010,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_10010);
		if (!D0 && !D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_00110,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_00110);
		if (!D0 && D2 && !D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_01010,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_01010);
		if (!D0 && D2 && D3 && S0 && !S1) (D1 +=> Z) = (`C12T32_LLUP0_MUX41X8_D1_R_Z_R_01110,`C12T32_LLUP0_MUX41X8_D1_F_Z_F_01110);
		if (!D0 && !D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_00001,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_00001);
		if (D0 && !D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_10101,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_10101);
		if (D0 && D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_11001,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_11001);
		if (D0 && D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_11101,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_11101);
		if (D0 && !D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_10001,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_10001);
		if (!D0 && !D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_00101,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_00101);
		if (!D0 && D1 && !D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_01001,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_01001);
		if (!D0 && D1 && D3 && !S0 && S1) (D2 +=> Z) = (`C12T32_LLUP0_MUX41X8_D2_R_Z_R_01101,`C12T32_LLUP0_MUX41X8_D2_F_Z_F_01101);
		if (!D0 && !D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_00011,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_00011);
		if (D0 && !D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_10111,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_10111);
		if (D0 && D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_11011,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_11011);
		if (D0 && D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_11111,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_11111);
		if (D0 && !D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_10011,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_10011);
		if (!D0 && !D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_00111,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_00111);
		if (!D0 && D1 && !D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_01011,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_01011);
		if (!D0 && D1 && D2 && S0 && S1) (D3 +=> Z) = (`C12T32_LLUP0_MUX41X8_D3_R_Z_R_01111,`C12T32_LLUP0_MUX41X8_D3_F_Z_F_01111);
		if (!D0 && !D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_00101,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_00101);
		if (D0 && !D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_10101,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_10101);
		if (D0 && !D1 && D2 && D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_10110,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_10110);
		if (D0 && D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_11101,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_11101);
		if (D0 && !D1 && D2 && !D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_10100,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_10100);
		if (!D0 && D1 && D2 && !D3 && S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_01101,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_01101);
		if (D0 && !D1 && !D2 && !D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_10000,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_10000);
		if (D0 && !D1 && !D2 && D3 && !S1) (S0 -=> Z) = (`C12T32_LLUP0_MUX41X8_S0_F_Z_R_10010,`C12T32_LLUP0_MUX41X8_S0_R_Z_F_10010);
		if (!D0 && !D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_00011,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_00011);
		if (!D0 && D1 && D2 && D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_01110,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_01110);
		if (D0 && !D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_10011,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_10011);
		if (D0 && D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_11011,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_11011);
		if (!D0 && D1 && D2 && !D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_01100,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_01100);
		if (!D0 && D1 && !D2 && !D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_01000,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_01000);
		if (!D0 && D1 && !D2 && D3 && !S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_01010,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_01010);
		if (!D0 && D1 && !D2 && D3 && S1) (S0 +=> Z) = (`C12T32_LLUP0_MUX41X8_S0_R_Z_R_01011,`C12T32_LLUP0_MUX41X8_S0_F_Z_F_01011);
		if (!D0 && D1 && !D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_01001,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_01001);
		if (D0 && D1 && !D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_11001,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_11001);
		if (D0 && D1 && !D2 && D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_11010,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_11010);
		if (D0 && D1 && D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_11101,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_11101);
		if (D0 && D1 && !D2 && !D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_11000,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_11000);
		if (!D0 && D1 && D2 && !D3 && S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_01101,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_01101);
		if (D0 && !D1 && !D2 && !D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_10000,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_10000);
		if (D0 && !D1 && !D2 && D3 && !S0) (S1 -=> Z) = (`C12T32_LLUP0_MUX41X8_S1_F_Z_R_10010,`C12T32_LLUP0_MUX41X8_S1_R_Z_F_10010);
		if (!D0 && !D1 && !D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_00011,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_00011);
		if (!D0 && D1 && D2 && D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_01110,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_01110);
		if (D0 && !D1 && !D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_10011,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_10011);
		if (D0 && !D1 && D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_10111,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_10111);
		if (!D0 && D1 && D2 && !D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_01100,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_01100);
		if (!D0 && !D1 && D2 && !D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_00100,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_00100);
		if (!D0 && !D1 && D2 && D3 && !S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_00110,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_00110);
		if (!D0 && !D1 && D2 && D3 && S0) (S1 +=> Z) = (`C12T32_LLUP0_MUX41X8_S1_R_Z_R_00111,`C12T32_LLUP0_MUX41X8_S1_F_Z_F_00111);


	endspecify

endmodule // C12T32_LLUP0_MUX41X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUXI21X10_D0_R_Z_F_00 0.1
`define C12T32_LLUP0_MUXI21X10_D0_F_Z_R_00 0.1
`define C12T32_LLUP0_MUXI21X10_D0_R_Z_F_10 0.1
`define C12T32_LLUP0_MUXI21X10_D0_F_Z_R_10 0.1
`define C12T32_LLUP0_MUXI21X10_D1_R_Z_F_01 0.1
`define C12T32_LLUP0_MUXI21X10_D1_F_Z_R_01 0.1
`define C12T32_LLUP0_MUXI21X10_D1_R_Z_F_11 0.1
`define C12T32_LLUP0_MUXI21X10_D1_F_Z_R_11 0.1
`define C12T32_LLUP0_MUXI21X10_S0_R_Z_F_01 0.1
`define C12T32_LLUP0_MUXI21X10_S0_F_Z_R_01 0.1
`define C12T32_LLUP0_MUXI21X10_S0_R_Z_R_10 0.1
`define C12T32_LLUP0_MUXI21X10_S0_F_Z_F_10 0.1

module C12T32_LLUP0_MUXI21X10 (Z, D0, D1, S0);

	output Z;
	input D0;
	input D1;
	input S0;

	U_MUX2   U1 (INTERNAL1, D0, D1, S0) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!D1 && !S0) (D0 -=> Z) = (`C12T32_LLUP0_MUXI21X10_D0_F_Z_R_00,`C12T32_LLUP0_MUXI21X10_D0_R_Z_F_00);
		if (D1 && !S0) (D0 -=> Z) = (`C12T32_LLUP0_MUXI21X10_D0_F_Z_R_10,`C12T32_LLUP0_MUXI21X10_D0_R_Z_F_10);
		if (!D0 && S0) (D1 -=> Z) = (`C12T32_LLUP0_MUXI21X10_D1_F_Z_R_01,`C12T32_LLUP0_MUXI21X10_D1_R_Z_F_01);
		if (D0 && S0) (D1 -=> Z) = (`C12T32_LLUP0_MUXI21X10_D1_F_Z_R_11,`C12T32_LLUP0_MUXI21X10_D1_R_Z_F_11);
		if (!D0 && D1) (S0 -=> Z) = (`C12T32_LLUP0_MUXI21X10_S0_F_Z_R_01,`C12T32_LLUP0_MUXI21X10_S0_R_Z_F_01);
		if (D0 && !D1) (S0 +=> Z) = (`C12T32_LLUP0_MUXI21X10_S0_R_Z_R_10,`C12T32_LLUP0_MUXI21X10_S0_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_MUXI21X10


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUXI21X21_D0_R_Z_F_00 0.1
`define C12T32_LLUP0_MUXI21X21_D0_F_Z_R_00 0.1
`define C12T32_LLUP0_MUXI21X21_D0_R_Z_F_10 0.1
`define C12T32_LLUP0_MUXI21X21_D0_F_Z_R_10 0.1
`define C12T32_LLUP0_MUXI21X21_D1_R_Z_F_01 0.1
`define C12T32_LLUP0_MUXI21X21_D1_F_Z_R_01 0.1
`define C12T32_LLUP0_MUXI21X21_D1_R_Z_F_11 0.1
`define C12T32_LLUP0_MUXI21X21_D1_F_Z_R_11 0.1
`define C12T32_LLUP0_MUXI21X21_S0_R_Z_F_01 0.1
`define C12T32_LLUP0_MUXI21X21_S0_F_Z_R_01 0.1
`define C12T32_LLUP0_MUXI21X21_S0_R_Z_R_10 0.1
`define C12T32_LLUP0_MUXI21X21_S0_F_Z_F_10 0.1

module C12T32_LLUP0_MUXI21X21 (Z, D0, D1, S0);

	output Z;
	input D0;
	input D1;
	input S0;

	U_MUX2   U1 (INTERNAL1, D0, D1, S0) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!D1 && !S0) (D0 -=> Z) = (`C12T32_LLUP0_MUXI21X21_D0_F_Z_R_00,`C12T32_LLUP0_MUXI21X21_D0_R_Z_F_00);
		if (D1 && !S0) (D0 -=> Z) = (`C12T32_LLUP0_MUXI21X21_D0_F_Z_R_10,`C12T32_LLUP0_MUXI21X21_D0_R_Z_F_10);
		if (!D0 && S0) (D1 -=> Z) = (`C12T32_LLUP0_MUXI21X21_D1_F_Z_R_01,`C12T32_LLUP0_MUXI21X21_D1_R_Z_F_01);
		if (D0 && S0) (D1 -=> Z) = (`C12T32_LLUP0_MUXI21X21_D1_F_Z_R_11,`C12T32_LLUP0_MUXI21X21_D1_R_Z_F_11);
		if (!D0 && D1) (S0 -=> Z) = (`C12T32_LLUP0_MUXI21X21_S0_F_Z_R_01,`C12T32_LLUP0_MUXI21X21_S0_R_Z_F_01);
		if (D0 && !D1) (S0 +=> Z) = (`C12T32_LLUP0_MUXI21X21_S0_R_Z_R_10,`C12T32_LLUP0_MUXI21X21_S0_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_MUXI21X21


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_MUXI21X5_D0_R_Z_F_00 0.1
`define C12T32_LLUP0_MUXI21X5_D0_F_Z_R_00 0.1
`define C12T32_LLUP0_MUXI21X5_D0_R_Z_F_10 0.1
`define C12T32_LLUP0_MUXI21X5_D0_F_Z_R_10 0.1
`define C12T32_LLUP0_MUXI21X5_D1_R_Z_F_01 0.1
`define C12T32_LLUP0_MUXI21X5_D1_F_Z_R_01 0.1
`define C12T32_LLUP0_MUXI21X5_D1_R_Z_F_11 0.1
`define C12T32_LLUP0_MUXI21X5_D1_F_Z_R_11 0.1
`define C12T32_LLUP0_MUXI21X5_S0_R_Z_F_01 0.1
`define C12T32_LLUP0_MUXI21X5_S0_F_Z_R_01 0.1
`define C12T32_LLUP0_MUXI21X5_S0_R_Z_R_10 0.1
`define C12T32_LLUP0_MUXI21X5_S0_F_Z_F_10 0.1

module C12T32_LLUP0_MUXI21X5 (Z, D0, D1, S0);

	output Z;
	input D0;
	input D1;
	input S0;

	U_MUX2   U1 (INTERNAL1, D0, D1, S0) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!D1 && !S0) (D0 -=> Z) = (`C12T32_LLUP0_MUXI21X5_D0_F_Z_R_00,`C12T32_LLUP0_MUXI21X5_D0_R_Z_F_00);
		if (D1 && !S0) (D0 -=> Z) = (`C12T32_LLUP0_MUXI21X5_D0_F_Z_R_10,`C12T32_LLUP0_MUXI21X5_D0_R_Z_F_10);
		if (!D0 && S0) (D1 -=> Z) = (`C12T32_LLUP0_MUXI21X5_D1_F_Z_R_01,`C12T32_LLUP0_MUXI21X5_D1_R_Z_F_01);
		if (D0 && S0) (D1 -=> Z) = (`C12T32_LLUP0_MUXI21X5_D1_F_Z_R_11,`C12T32_LLUP0_MUXI21X5_D1_R_Z_F_11);
		if (!D0 && D1) (S0 -=> Z) = (`C12T32_LLUP0_MUXI21X5_S0_F_Z_R_01,`C12T32_LLUP0_MUXI21X5_S0_R_Z_F_01);
		if (D0 && !D1) (S0 +=> Z) = (`C12T32_LLUP0_MUXI21X5_S0_R_Z_R_10,`C12T32_LLUP0_MUXI21X5_S0_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_MUXI21X5


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X11_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X11_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X11_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X11_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X11 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X11_A_F_Z_R_1,`C12T32_LLUP0_NAND2X11_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X11_B_F_Z_R_1,`C12T32_LLUP0_NAND2X11_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X11


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X13_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X13_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X13_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X13_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X13 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X13_A_F_Z_R_1,`C12T32_LLUP0_NAND2X13_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X13_B_F_Z_R_1,`C12T32_LLUP0_NAND2X13_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X13


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X20_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X20_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X20_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X20_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X20 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X20_A_F_Z_R_1,`C12T32_LLUP0_NAND2X20_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X20_B_F_Z_R_1,`C12T32_LLUP0_NAND2X20_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X20


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X22_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X22_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X22_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X22_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X22 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X22_A_F_Z_R_1,`C12T32_LLUP0_NAND2X22_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X22_B_F_Z_R_1,`C12T32_LLUP0_NAND2X22_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X22


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X3_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X3_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X3_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X3_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X3 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X3_A_F_Z_R_1,`C12T32_LLUP0_NAND2X3_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X3_B_F_Z_R_1,`C12T32_LLUP0_NAND2X3_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X3


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X5_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X5_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X5_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X5_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X5 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X5_A_F_Z_R_1,`C12T32_LLUP0_NAND2X5_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X5_B_F_Z_R_1,`C12T32_LLUP0_NAND2X5_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X5


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND2X7_A_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X7_A_F_Z_R_1 0.1
`define C12T32_LLUP0_NAND2X7_B_R_Z_F_1 0.1
`define C12T32_LLUP0_NAND2X7_B_F_Z_R_1 0.1

module C12T32_LLUP0_NAND2X7 (Z, A, B);

	output Z;
	input A;
	input B;

	and    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A -=> Z) = (`C12T32_LLUP0_NAND2X7_A_F_Z_R_1,`C12T32_LLUP0_NAND2X7_A_R_Z_F_1);
		if (A) (B -=> Z) = (`C12T32_LLUP0_NAND2X7_B_F_Z_R_1,`C12T32_LLUP0_NAND2X7_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_NAND2X7


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND3X12_A_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X12_A_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X12_B_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X12_B_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X12_C_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X12_C_F_Z_R_11 0.1

module C12T32_LLUP0_NAND3X12 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_NAND3X12_A_F_Z_R_11,`C12T32_LLUP0_NAND3X12_A_R_Z_F_11);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_NAND3X12_B_F_Z_R_11,`C12T32_LLUP0_NAND3X12_B_R_Z_F_11);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_NAND3X12_C_F_Z_R_11,`C12T32_LLUP0_NAND3X12_C_R_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_NAND3X12


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND3X15_A_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X15_A_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X15_B_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X15_B_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X15_C_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X15_C_F_Z_R_11 0.1

module C12T32_LLUP0_NAND3X15 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_NAND3X15_A_F_Z_R_11,`C12T32_LLUP0_NAND3X15_A_R_Z_F_11);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_NAND3X15_B_F_Z_R_11,`C12T32_LLUP0_NAND3X15_B_R_Z_F_11);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_NAND3X15_C_F_Z_R_11,`C12T32_LLUP0_NAND3X15_C_R_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_NAND3X15


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND3X18_A_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X18_A_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X18_B_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X18_B_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X18_C_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X18_C_F_Z_R_11 0.1

module C12T32_LLUP0_NAND3X18 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_NAND3X18_A_F_Z_R_11,`C12T32_LLUP0_NAND3X18_A_R_Z_F_11);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_NAND3X18_B_F_Z_R_11,`C12T32_LLUP0_NAND3X18_B_R_Z_F_11);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_NAND3X18_C_F_Z_R_11,`C12T32_LLUP0_NAND3X18_C_R_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_NAND3X18


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND3X4_A_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X4_A_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X4_B_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X4_B_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X4_C_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X4_C_F_Z_R_11 0.1

module C12T32_LLUP0_NAND3X4 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_NAND3X4_A_F_Z_R_11,`C12T32_LLUP0_NAND3X4_A_R_Z_F_11);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_NAND3X4_B_F_Z_R_11,`C12T32_LLUP0_NAND3X4_B_R_Z_F_11);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_NAND3X4_C_F_Z_R_11,`C12T32_LLUP0_NAND3X4_C_R_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_NAND3X4


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND3X6_A_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X6_A_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X6_B_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X6_B_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X6_C_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X6_C_F_Z_R_11 0.1

module C12T32_LLUP0_NAND3X6 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_NAND3X6_A_F_Z_R_11,`C12T32_LLUP0_NAND3X6_A_R_Z_F_11);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_NAND3X6_B_F_Z_R_11,`C12T32_LLUP0_NAND3X6_B_R_Z_F_11);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_NAND3X6_C_F_Z_R_11,`C12T32_LLUP0_NAND3X6_C_R_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_NAND3X6


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NAND3X7_A_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X7_A_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X7_B_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X7_B_F_Z_R_11 0.1
`define C12T32_LLUP0_NAND3X7_C_R_Z_F_11 0.1
`define C12T32_LLUP0_NAND3X7_C_F_Z_R_11 0.1

module C12T32_LLUP0_NAND3X7 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	and    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_NAND3X7_A_F_Z_R_11,`C12T32_LLUP0_NAND3X7_A_R_Z_F_11);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_NAND3X7_B_F_Z_R_11,`C12T32_LLUP0_NAND3X7_B_R_Z_F_11);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_NAND3X7_C_F_Z_R_11,`C12T32_LLUP0_NAND3X7_C_R_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_NAND3X7


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X11_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X11_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X11_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X11_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X11 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X11_A_F_Z_R_0,`C12T32_LLUP0_NOR2X11_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X11_B_F_Z_R_0,`C12T32_LLUP0_NOR2X11_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X11


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X14_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X14_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X14_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X14_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X14 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X14_A_F_Z_R_0,`C12T32_LLUP0_NOR2X14_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X14_B_F_Z_R_0,`C12T32_LLUP0_NOR2X14_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X14


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X21_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X21_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X21_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X21_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X21 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X21_A_F_Z_R_0,`C12T32_LLUP0_NOR2X21_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X21_B_F_Z_R_0,`C12T32_LLUP0_NOR2X21_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X21


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X22_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X22_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X22_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X22_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X22 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X22_A_F_Z_R_0,`C12T32_LLUP0_NOR2X22_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X22_B_F_Z_R_0,`C12T32_LLUP0_NOR2X22_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X22


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X3_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X3_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X3_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X3_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X3 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X3_A_F_Z_R_0,`C12T32_LLUP0_NOR2X3_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X3_B_F_Z_R_0,`C12T32_LLUP0_NOR2X3_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X3


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X5_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X5_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X5_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X5_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X5 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X5_A_F_Z_R_0,`C12T32_LLUP0_NOR2X5_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X5_B_F_Z_R_0,`C12T32_LLUP0_NOR2X5_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X5


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR2X7_A_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X7_A_F_Z_R_0 0.1
`define C12T32_LLUP0_NOR2X7_B_R_Z_F_0 0.1
`define C12T32_LLUP0_NOR2X7_B_F_Z_R_0 0.1

module C12T32_LLUP0_NOR2X7 (Z, A, B);

	output Z;
	input A;
	input B;

	or    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B) (A -=> Z) = (`C12T32_LLUP0_NOR2X7_A_F_Z_R_0,`C12T32_LLUP0_NOR2X7_A_R_Z_F_0);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_NOR2X7_B_F_Z_R_0,`C12T32_LLUP0_NOR2X7_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_NOR2X7


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR3X13_A_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X13_A_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X13_B_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X13_B_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X13_C_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X13_C_F_Z_R_00 0.1

module C12T32_LLUP0_NOR3X13 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_NOR3X13_A_F_Z_R_00,`C12T32_LLUP0_NOR3X13_A_R_Z_F_00);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_NOR3X13_B_F_Z_R_00,`C12T32_LLUP0_NOR3X13_B_R_Z_F_00);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_NOR3X13_C_F_Z_R_00,`C12T32_LLUP0_NOR3X13_C_R_Z_F_00);


	endspecify

endmodule // C12T32_LLUP0_NOR3X13


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR3X15_A_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X15_A_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X15_B_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X15_B_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X15_C_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X15_C_F_Z_R_00 0.1

module C12T32_LLUP0_NOR3X15 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_NOR3X15_A_F_Z_R_00,`C12T32_LLUP0_NOR3X15_A_R_Z_F_00);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_NOR3X15_B_F_Z_R_00,`C12T32_LLUP0_NOR3X15_B_R_Z_F_00);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_NOR3X15_C_F_Z_R_00,`C12T32_LLUP0_NOR3X15_C_R_Z_F_00);


	endspecify

endmodule // C12T32_LLUP0_NOR3X15


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR3X19_A_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X19_A_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X19_B_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X19_B_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X19_C_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X19_C_F_Z_R_00 0.1

module C12T32_LLUP0_NOR3X19 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_NOR3X19_A_F_Z_R_00,`C12T32_LLUP0_NOR3X19_A_R_Z_F_00);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_NOR3X19_B_F_Z_R_00,`C12T32_LLUP0_NOR3X19_B_R_Z_F_00);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_NOR3X19_C_F_Z_R_00,`C12T32_LLUP0_NOR3X19_C_R_Z_F_00);


	endspecify

endmodule // C12T32_LLUP0_NOR3X19


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR3X4_A_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X4_A_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X4_B_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X4_B_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X4_C_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X4_C_F_Z_R_00 0.1

module C12T32_LLUP0_NOR3X4 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_NOR3X4_A_F_Z_R_00,`C12T32_LLUP0_NOR3X4_A_R_Z_F_00);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_NOR3X4_B_F_Z_R_00,`C12T32_LLUP0_NOR3X4_B_R_Z_F_00);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_NOR3X4_C_F_Z_R_00,`C12T32_LLUP0_NOR3X4_C_R_Z_F_00);


	endspecify

endmodule // C12T32_LLUP0_NOR3X4


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR3X6_A_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X6_A_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X6_B_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X6_B_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X6_C_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X6_C_F_Z_R_00 0.1

module C12T32_LLUP0_NOR3X6 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_NOR3X6_A_F_Z_R_00,`C12T32_LLUP0_NOR3X6_A_R_Z_F_00);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_NOR3X6_B_F_Z_R_00,`C12T32_LLUP0_NOR3X6_B_R_Z_F_00);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_NOR3X6_C_F_Z_R_00,`C12T32_LLUP0_NOR3X6_C_R_Z_F_00);


	endspecify

endmodule // C12T32_LLUP0_NOR3X6


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_NOR3X8_A_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X8_A_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X8_B_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X8_B_F_Z_R_00 0.1
`define C12T32_LLUP0_NOR3X8_C_R_Z_F_00 0.1
`define C12T32_LLUP0_NOR3X8_C_F_Z_R_00 0.1

module C12T32_LLUP0_NOR3X8 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_NOR3X8_A_F_Z_R_00,`C12T32_LLUP0_NOR3X8_A_R_Z_F_00);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_NOR3X8_B_F_Z_R_00,`C12T32_LLUP0_NOR3X8_B_R_Z_F_00);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_NOR3X8_C_F_Z_R_00,`C12T32_LLUP0_NOR3X8_C_R_Z_F_00);


	endspecify

endmodule // C12T32_LLUP0_NOR3X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA112X17_A_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X17_A_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X17_B_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X17_B_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X17_C_R_Z_R_101 0.1
`define C12T32_LLUP0_OA112X17_C_F_Z_F_101 0.1
`define C12T32_LLUP0_OA112X17_C_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X17_C_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X17_C_R_Z_R_111 0.1
`define C12T32_LLUP0_OA112X17_C_F_Z_F_111 0.1
`define C12T32_LLUP0_OA112X17_D_R_Z_R_101 0.1
`define C12T32_LLUP0_OA112X17_D_F_Z_F_101 0.1
`define C12T32_LLUP0_OA112X17_D_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X17_D_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X17_D_R_Z_R_111 0.1
`define C12T32_LLUP0_OA112X17_D_F_Z_F_111 0.1

module C12T32_LLUP0_OA112X17 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	or    U1 (INTERNAL1, A, B) ;
	and   #1 U2 (Z, INTERNAL1, C, D) ;



	specify

		if (!B && C && D) (A +=> Z) = (`C12T32_LLUP0_OA112X17_A_R_Z_R_011,`C12T32_LLUP0_OA112X17_A_F_Z_F_011);
		if (!A && C && D) (B +=> Z) = (`C12T32_LLUP0_OA112X17_B_R_Z_R_011,`C12T32_LLUP0_OA112X17_B_F_Z_F_011);
		if (A && !B && D) (C +=> Z) = (`C12T32_LLUP0_OA112X17_C_R_Z_R_101,`C12T32_LLUP0_OA112X17_C_F_Z_F_101);
		if (!A && B && D) (C +=> Z) = (`C12T32_LLUP0_OA112X17_C_R_Z_R_011,`C12T32_LLUP0_OA112X17_C_F_Z_F_011);
		if (A && B && D) (C +=> Z) = (`C12T32_LLUP0_OA112X17_C_R_Z_R_111,`C12T32_LLUP0_OA112X17_C_F_Z_F_111);
		if (A && !B && C) (D +=> Z) = (`C12T32_LLUP0_OA112X17_D_R_Z_R_101,`C12T32_LLUP0_OA112X17_D_F_Z_F_101);
		if (!A && B && C) (D +=> Z) = (`C12T32_LLUP0_OA112X17_D_R_Z_R_011,`C12T32_LLUP0_OA112X17_D_F_Z_F_011);
		if (A && B && C) (D +=> Z) = (`C12T32_LLUP0_OA112X17_D_R_Z_R_111,`C12T32_LLUP0_OA112X17_D_F_Z_F_111);


	endspecify

endmodule // C12T32_LLUP0_OA112X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA112X8_A_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X8_A_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X8_B_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X8_B_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X8_C_R_Z_R_101 0.1
`define C12T32_LLUP0_OA112X8_C_F_Z_F_101 0.1
`define C12T32_LLUP0_OA112X8_C_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X8_C_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X8_C_R_Z_R_111 0.1
`define C12T32_LLUP0_OA112X8_C_F_Z_F_111 0.1
`define C12T32_LLUP0_OA112X8_D_R_Z_R_101 0.1
`define C12T32_LLUP0_OA112X8_D_F_Z_F_101 0.1
`define C12T32_LLUP0_OA112X8_D_R_Z_R_011 0.1
`define C12T32_LLUP0_OA112X8_D_F_Z_F_011 0.1
`define C12T32_LLUP0_OA112X8_D_R_Z_R_111 0.1
`define C12T32_LLUP0_OA112X8_D_F_Z_F_111 0.1

module C12T32_LLUP0_OA112X8 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	or    U1 (INTERNAL1, A, B) ;
	and   #1 U2 (Z, INTERNAL1, C, D) ;



	specify

		if (!B && C && D) (A +=> Z) = (`C12T32_LLUP0_OA112X8_A_R_Z_R_011,`C12T32_LLUP0_OA112X8_A_F_Z_F_011);
		if (!A && C && D) (B +=> Z) = (`C12T32_LLUP0_OA112X8_B_R_Z_R_011,`C12T32_LLUP0_OA112X8_B_F_Z_F_011);
		if (A && !B && D) (C +=> Z) = (`C12T32_LLUP0_OA112X8_C_R_Z_R_101,`C12T32_LLUP0_OA112X8_C_F_Z_F_101);
		if (!A && B && D) (C +=> Z) = (`C12T32_LLUP0_OA112X8_C_R_Z_R_011,`C12T32_LLUP0_OA112X8_C_F_Z_F_011);
		if (A && B && D) (C +=> Z) = (`C12T32_LLUP0_OA112X8_C_R_Z_R_111,`C12T32_LLUP0_OA112X8_C_F_Z_F_111);
		if (A && !B && C) (D +=> Z) = (`C12T32_LLUP0_OA112X8_D_R_Z_R_101,`C12T32_LLUP0_OA112X8_D_F_Z_F_101);
		if (!A && B && C) (D +=> Z) = (`C12T32_LLUP0_OA112X8_D_R_Z_R_011,`C12T32_LLUP0_OA112X8_D_F_Z_F_011);
		if (A && B && C) (D +=> Z) = (`C12T32_LLUP0_OA112X8_D_R_Z_R_111,`C12T32_LLUP0_OA112X8_D_F_Z_F_111);


	endspecify

endmodule // C12T32_LLUP0_OA112X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA12X17_A_R_Z_R_01 0.1
`define C12T32_LLUP0_OA12X17_A_F_Z_F_01 0.1
`define C12T32_LLUP0_OA12X17_B_R_Z_R_01 0.1
`define C12T32_LLUP0_OA12X17_B_F_Z_F_01 0.1
`define C12T32_LLUP0_OA12X17_C_R_Z_R_01 0.1
`define C12T32_LLUP0_OA12X17_C_F_Z_F_01 0.1
`define C12T32_LLUP0_OA12X17_C_R_Z_R_11 0.1
`define C12T32_LLUP0_OA12X17_C_F_Z_F_11 0.1
`define C12T32_LLUP0_OA12X17_C_R_Z_R_10 0.1
`define C12T32_LLUP0_OA12X17_C_F_Z_F_10 0.1

module C12T32_LLUP0_OA12X17 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B) ;
	and   #1 U2 (Z, INTERNAL1, C) ;



	specify

		if (!B && C) (A +=> Z) = (`C12T32_LLUP0_OA12X17_A_R_Z_R_01,`C12T32_LLUP0_OA12X17_A_F_Z_F_01);
		if (!A && C) (B +=> Z) = (`C12T32_LLUP0_OA12X17_B_R_Z_R_01,`C12T32_LLUP0_OA12X17_B_F_Z_F_01);
		if (!A && B) (C +=> Z) = (`C12T32_LLUP0_OA12X17_C_R_Z_R_01,`C12T32_LLUP0_OA12X17_C_F_Z_F_01);
		if (A && B) (C +=> Z) = (`C12T32_LLUP0_OA12X17_C_R_Z_R_11,`C12T32_LLUP0_OA12X17_C_F_Z_F_11);
		if (A && !B) (C +=> Z) = (`C12T32_LLUP0_OA12X17_C_R_Z_R_10,`C12T32_LLUP0_OA12X17_C_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_OA12X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA12X8_A_R_Z_R_01 0.1
`define C12T32_LLUP0_OA12X8_A_F_Z_F_01 0.1
`define C12T32_LLUP0_OA12X8_B_R_Z_R_01 0.1
`define C12T32_LLUP0_OA12X8_B_F_Z_F_01 0.1
`define C12T32_LLUP0_OA12X8_C_R_Z_R_01 0.1
`define C12T32_LLUP0_OA12X8_C_F_Z_F_01 0.1
`define C12T32_LLUP0_OA12X8_C_R_Z_R_11 0.1
`define C12T32_LLUP0_OA12X8_C_F_Z_F_11 0.1
`define C12T32_LLUP0_OA12X8_C_R_Z_R_10 0.1
`define C12T32_LLUP0_OA12X8_C_F_Z_F_10 0.1

module C12T32_LLUP0_OA12X8 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL1, A, B) ;
	and   #1 U2 (Z, INTERNAL1, C) ;



	specify

		if (!B && C) (A +=> Z) = (`C12T32_LLUP0_OA12X8_A_R_Z_R_01,`C12T32_LLUP0_OA12X8_A_F_Z_F_01);
		if (!A && C) (B +=> Z) = (`C12T32_LLUP0_OA12X8_B_R_Z_R_01,`C12T32_LLUP0_OA12X8_B_F_Z_F_01);
		if (!A && B) (C +=> Z) = (`C12T32_LLUP0_OA12X8_C_R_Z_R_01,`C12T32_LLUP0_OA12X8_C_F_Z_F_01);
		if (A && B) (C +=> Z) = (`C12T32_LLUP0_OA12X8_C_R_Z_R_11,`C12T32_LLUP0_OA12X8_C_F_Z_F_11);
		if (A && !B) (C +=> Z) = (`C12T32_LLUP0_OA12X8_C_R_Z_R_10,`C12T32_LLUP0_OA12X8_C_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_OA12X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA222X17_A_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_01110 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_01111 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_01111 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_01101 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_01101 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_00110 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_00110 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_00101 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_00101 0.1
`define C12T32_LLUP0_OA222X17_A_R_Z_R_00111 0.1
`define C12T32_LLUP0_OA222X17_A_F_Z_F_00111 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_01110 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_01111 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_01111 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_01101 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_01101 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_00110 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_00110 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_00101 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_00101 0.1
`define C12T32_LLUP0_OA222X17_B_R_Z_R_00111 0.1
`define C12T32_LLUP0_OA222X17_B_F_Z_F_00111 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_11011 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_11011 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_10001 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_10001 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_10011 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_10011 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_11001 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_11001 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X17_C_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X17_C_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_11011 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_11011 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_10001 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_10001 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_10011 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_10011 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_11001 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_11001 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X17_D_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X17_D_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_11100 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_11100 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_11110 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_11110 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_10110 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_10110 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_10100 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_10100 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_01100 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_01100 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X17_E_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X17_E_F_Z_F_01110 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_11100 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_11100 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_11110 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_11110 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_10110 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_10110 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_10100 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_10100 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_01100 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_01100 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X17_F_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X17_F_F_Z_F_01110 0.1

module C12T32_LLUP0_OA222X17 (Z, A, B, C, D, E, F);

	output Z;
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;

	or    U1 (INTERNAL2, A, B) ;
	or    U2 (INTERNAL3, C, D) ;
	or    U3 (INTERNAL4, E, F) ;
	and    U4 (INTERNAL1, INTERNAL2, INTERNAL3, INTERNAL4) ;
	not    U5 (NET1, INTERNAL1) ;
	not   #1 U6 (Z, NET1) ;



	specify

		if (!B && C && D && E && !F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_01110,`C12T32_LLUP0_OA222X17_A_F_Z_F_01110);
		if (!B && C && D && E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_01111,`C12T32_LLUP0_OA222X17_A_F_Z_F_01111);
		if (!B && C && !D && !E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_01001,`C12T32_LLUP0_OA222X17_A_F_Z_F_01001);
		if (!B && C && !D && E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_01011,`C12T32_LLUP0_OA222X17_A_F_Z_F_01011);
		if (!B && C && !D && E && !F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_01010,`C12T32_LLUP0_OA222X17_A_F_Z_F_01010);
		if (!B && C && D && !E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_01101,`C12T32_LLUP0_OA222X17_A_F_Z_F_01101);
		if (!B && !C && D && E && !F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_00110,`C12T32_LLUP0_OA222X17_A_F_Z_F_00110);
		if (!B && !C && D && !E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_00101,`C12T32_LLUP0_OA222X17_A_F_Z_F_00101);
		if (!B && !C && D && E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X17_A_R_Z_R_00111,`C12T32_LLUP0_OA222X17_A_F_Z_F_00111);
		if (!A && C && D && E && !F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_01110,`C12T32_LLUP0_OA222X17_B_F_Z_F_01110);
		if (!A && C && D && E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_01111,`C12T32_LLUP0_OA222X17_B_F_Z_F_01111);
		if (!A && C && !D && !E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_01001,`C12T32_LLUP0_OA222X17_B_F_Z_F_01001);
		if (!A && C && !D && E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_01011,`C12T32_LLUP0_OA222X17_B_F_Z_F_01011);
		if (!A && C && !D && E && !F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_01010,`C12T32_LLUP0_OA222X17_B_F_Z_F_01010);
		if (!A && C && D && !E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_01101,`C12T32_LLUP0_OA222X17_B_F_Z_F_01101);
		if (!A && !C && D && E && !F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_00110,`C12T32_LLUP0_OA222X17_B_F_Z_F_00110);
		if (!A && !C && D && !E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_00101,`C12T32_LLUP0_OA222X17_B_F_Z_F_00101);
		if (!A && !C && D && E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X17_B_R_Z_R_00111,`C12T32_LLUP0_OA222X17_B_F_Z_F_00111);
		if (A && B && !D && E && !F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_11010,`C12T32_LLUP0_OA222X17_C_F_Z_F_11010);
		if (A && B && !D && E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_11011,`C12T32_LLUP0_OA222X17_C_F_Z_F_11011);
		if (A && !B && !D && !E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_10001,`C12T32_LLUP0_OA222X17_C_F_Z_F_10001);
		if (A && !B && !D && E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_10011,`C12T32_LLUP0_OA222X17_C_F_Z_F_10011);
		if (A && !B && !D && E && !F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_10010,`C12T32_LLUP0_OA222X17_C_F_Z_F_10010);
		if (A && B && !D && !E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_11001,`C12T32_LLUP0_OA222X17_C_F_Z_F_11001);
		if (!A && B && !D && E && !F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_01010,`C12T32_LLUP0_OA222X17_C_F_Z_F_01010);
		if (!A && B && !D && !E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_01001,`C12T32_LLUP0_OA222X17_C_F_Z_F_01001);
		if (!A && B && !D && E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X17_C_R_Z_R_01011,`C12T32_LLUP0_OA222X17_C_F_Z_F_01011);
		if (A && B && !C && E && !F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_11010,`C12T32_LLUP0_OA222X17_D_F_Z_F_11010);
		if (A && B && !C && E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_11011,`C12T32_LLUP0_OA222X17_D_F_Z_F_11011);
		if (A && !B && !C && !E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_10001,`C12T32_LLUP0_OA222X17_D_F_Z_F_10001);
		if (A && !B && !C && E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_10011,`C12T32_LLUP0_OA222X17_D_F_Z_F_10011);
		if (A && !B && !C && E && !F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_10010,`C12T32_LLUP0_OA222X17_D_F_Z_F_10010);
		if (A && B && !C && !E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_11001,`C12T32_LLUP0_OA222X17_D_F_Z_F_11001);
		if (!A && B && !C && E && !F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_01010,`C12T32_LLUP0_OA222X17_D_F_Z_F_01010);
		if (!A && B && !C && !E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_01001,`C12T32_LLUP0_OA222X17_D_F_Z_F_01001);
		if (!A && B && !C && E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X17_D_R_Z_R_01011,`C12T32_LLUP0_OA222X17_D_F_Z_F_01011);
		if (A && B && C && !D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_11100,`C12T32_LLUP0_OA222X17_E_F_Z_F_11100);
		if (A && B && C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_11110,`C12T32_LLUP0_OA222X17_E_F_Z_F_11110);
		if (A && !B && !C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_10010,`C12T32_LLUP0_OA222X17_E_F_Z_F_10010);
		if (A && !B && C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_10110,`C12T32_LLUP0_OA222X17_E_F_Z_F_10110);
		if (A && !B && C && !D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_10100,`C12T32_LLUP0_OA222X17_E_F_Z_F_10100);
		if (A && B && !C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_11010,`C12T32_LLUP0_OA222X17_E_F_Z_F_11010);
		if (!A && B && C && !D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_01100,`C12T32_LLUP0_OA222X17_E_F_Z_F_01100);
		if (!A && B && !C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_01010,`C12T32_LLUP0_OA222X17_E_F_Z_F_01010);
		if (!A && B && C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X17_E_R_Z_R_01110,`C12T32_LLUP0_OA222X17_E_F_Z_F_01110);
		if (A && B && C && !D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_11100,`C12T32_LLUP0_OA222X17_F_F_Z_F_11100);
		if (A && B && C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_11110,`C12T32_LLUP0_OA222X17_F_F_Z_F_11110);
		if (A && !B && !C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_10010,`C12T32_LLUP0_OA222X17_F_F_Z_F_10010);
		if (A && !B && C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_10110,`C12T32_LLUP0_OA222X17_F_F_Z_F_10110);
		if (A && !B && C && !D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_10100,`C12T32_LLUP0_OA222X17_F_F_Z_F_10100);
		if (A && B && !C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_11010,`C12T32_LLUP0_OA222X17_F_F_Z_F_11010);
		if (!A && B && C && !D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_01100,`C12T32_LLUP0_OA222X17_F_F_Z_F_01100);
		if (!A && B && !C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_01010,`C12T32_LLUP0_OA222X17_F_F_Z_F_01010);
		if (!A && B && C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X17_F_R_Z_R_01110,`C12T32_LLUP0_OA222X17_F_F_Z_F_01110);


	endspecify

endmodule // C12T32_LLUP0_OA222X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA222X8_A_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_01110 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_01111 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_01111 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_01101 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_01101 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_00110 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_00110 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_00101 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_00101 0.1
`define C12T32_LLUP0_OA222X8_A_R_Z_R_00111 0.1
`define C12T32_LLUP0_OA222X8_A_F_Z_F_00111 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_01110 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_01111 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_01111 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_01101 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_01101 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_00110 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_00110 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_00101 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_00101 0.1
`define C12T32_LLUP0_OA222X8_B_R_Z_R_00111 0.1
`define C12T32_LLUP0_OA222X8_B_F_Z_F_00111 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_11011 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_11011 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_10001 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_10001 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_10011 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_10011 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_11001 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_11001 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X8_C_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X8_C_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_11011 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_11011 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_10001 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_10001 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_10011 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_10011 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_11001 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_11001 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_01001 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_01001 0.1
`define C12T32_LLUP0_OA222X8_D_R_Z_R_01011 0.1
`define C12T32_LLUP0_OA222X8_D_F_Z_F_01011 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_11100 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_11100 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_11110 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_11110 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_10110 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_10110 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_10100 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_10100 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_01100 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_01100 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X8_E_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X8_E_F_Z_F_01110 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_11100 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_11100 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_11110 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_11110 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_10010 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_10010 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_10110 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_10110 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_10100 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_10100 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_11010 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_11010 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_01100 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_01100 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_01010 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_01010 0.1
`define C12T32_LLUP0_OA222X8_F_R_Z_R_01110 0.1
`define C12T32_LLUP0_OA222X8_F_F_Z_F_01110 0.1

module C12T32_LLUP0_OA222X8 (Z, A, B, C, D, E, F);

	output Z;
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;

	or    U1 (INTERNAL2, A, B) ;
	or    U2 (INTERNAL3, C, D) ;
	or    U3 (INTERNAL4, E, F) ;
	and    U4 (INTERNAL1, INTERNAL2, INTERNAL3, INTERNAL4) ;
	not    U5 (NET1, INTERNAL1) ;
	not   #1 U6 (Z, NET1) ;



	specify

		if (!B && C && D && E && !F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_01110,`C12T32_LLUP0_OA222X8_A_F_Z_F_01110);
		if (!B && C && D && E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_01111,`C12T32_LLUP0_OA222X8_A_F_Z_F_01111);
		if (!B && C && !D && !E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_01001,`C12T32_LLUP0_OA222X8_A_F_Z_F_01001);
		if (!B && C && !D && E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_01011,`C12T32_LLUP0_OA222X8_A_F_Z_F_01011);
		if (!B && C && !D && E && !F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_01010,`C12T32_LLUP0_OA222X8_A_F_Z_F_01010);
		if (!B && C && D && !E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_01101,`C12T32_LLUP0_OA222X8_A_F_Z_F_01101);
		if (!B && !C && D && E && !F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_00110,`C12T32_LLUP0_OA222X8_A_F_Z_F_00110);
		if (!B && !C && D && !E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_00101,`C12T32_LLUP0_OA222X8_A_F_Z_F_00101);
		if (!B && !C && D && E && F) (A +=> Z) = (`C12T32_LLUP0_OA222X8_A_R_Z_R_00111,`C12T32_LLUP0_OA222X8_A_F_Z_F_00111);
		if (!A && C && D && E && !F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_01110,`C12T32_LLUP0_OA222X8_B_F_Z_F_01110);
		if (!A && C && D && E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_01111,`C12T32_LLUP0_OA222X8_B_F_Z_F_01111);
		if (!A && C && !D && !E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_01001,`C12T32_LLUP0_OA222X8_B_F_Z_F_01001);
		if (!A && C && !D && E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_01011,`C12T32_LLUP0_OA222X8_B_F_Z_F_01011);
		if (!A && C && !D && E && !F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_01010,`C12T32_LLUP0_OA222X8_B_F_Z_F_01010);
		if (!A && C && D && !E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_01101,`C12T32_LLUP0_OA222X8_B_F_Z_F_01101);
		if (!A && !C && D && E && !F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_00110,`C12T32_LLUP0_OA222X8_B_F_Z_F_00110);
		if (!A && !C && D && !E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_00101,`C12T32_LLUP0_OA222X8_B_F_Z_F_00101);
		if (!A && !C && D && E && F) (B +=> Z) = (`C12T32_LLUP0_OA222X8_B_R_Z_R_00111,`C12T32_LLUP0_OA222X8_B_F_Z_F_00111);
		if (A && B && !D && E && !F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_11010,`C12T32_LLUP0_OA222X8_C_F_Z_F_11010);
		if (A && B && !D && E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_11011,`C12T32_LLUP0_OA222X8_C_F_Z_F_11011);
		if (A && !B && !D && !E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_10001,`C12T32_LLUP0_OA222X8_C_F_Z_F_10001);
		if (A && !B && !D && E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_10011,`C12T32_LLUP0_OA222X8_C_F_Z_F_10011);
		if (A && !B && !D && E && !F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_10010,`C12T32_LLUP0_OA222X8_C_F_Z_F_10010);
		if (A && B && !D && !E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_11001,`C12T32_LLUP0_OA222X8_C_F_Z_F_11001);
		if (!A && B && !D && E && !F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_01010,`C12T32_LLUP0_OA222X8_C_F_Z_F_01010);
		if (!A && B && !D && !E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_01001,`C12T32_LLUP0_OA222X8_C_F_Z_F_01001);
		if (!A && B && !D && E && F) (C +=> Z) = (`C12T32_LLUP0_OA222X8_C_R_Z_R_01011,`C12T32_LLUP0_OA222X8_C_F_Z_F_01011);
		if (A && B && !C && E && !F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_11010,`C12T32_LLUP0_OA222X8_D_F_Z_F_11010);
		if (A && B && !C && E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_11011,`C12T32_LLUP0_OA222X8_D_F_Z_F_11011);
		if (A && !B && !C && !E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_10001,`C12T32_LLUP0_OA222X8_D_F_Z_F_10001);
		if (A && !B && !C && E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_10011,`C12T32_LLUP0_OA222X8_D_F_Z_F_10011);
		if (A && !B && !C && E && !F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_10010,`C12T32_LLUP0_OA222X8_D_F_Z_F_10010);
		if (A && B && !C && !E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_11001,`C12T32_LLUP0_OA222X8_D_F_Z_F_11001);
		if (!A && B && !C && E && !F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_01010,`C12T32_LLUP0_OA222X8_D_F_Z_F_01010);
		if (!A && B && !C && !E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_01001,`C12T32_LLUP0_OA222X8_D_F_Z_F_01001);
		if (!A && B && !C && E && F) (D +=> Z) = (`C12T32_LLUP0_OA222X8_D_R_Z_R_01011,`C12T32_LLUP0_OA222X8_D_F_Z_F_01011);
		if (A && B && C && !D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_11100,`C12T32_LLUP0_OA222X8_E_F_Z_F_11100);
		if (A && B && C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_11110,`C12T32_LLUP0_OA222X8_E_F_Z_F_11110);
		if (A && !B && !C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_10010,`C12T32_LLUP0_OA222X8_E_F_Z_F_10010);
		if (A && !B && C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_10110,`C12T32_LLUP0_OA222X8_E_F_Z_F_10110);
		if (A && !B && C && !D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_10100,`C12T32_LLUP0_OA222X8_E_F_Z_F_10100);
		if (A && B && !C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_11010,`C12T32_LLUP0_OA222X8_E_F_Z_F_11010);
		if (!A && B && C && !D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_01100,`C12T32_LLUP0_OA222X8_E_F_Z_F_01100);
		if (!A && B && !C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_01010,`C12T32_LLUP0_OA222X8_E_F_Z_F_01010);
		if (!A && B && C && D && !F) (E +=> Z) = (`C12T32_LLUP0_OA222X8_E_R_Z_R_01110,`C12T32_LLUP0_OA222X8_E_F_Z_F_01110);
		if (A && B && C && !D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_11100,`C12T32_LLUP0_OA222X8_F_F_Z_F_11100);
		if (A && B && C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_11110,`C12T32_LLUP0_OA222X8_F_F_Z_F_11110);
		if (A && !B && !C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_10010,`C12T32_LLUP0_OA222X8_F_F_Z_F_10010);
		if (A && !B && C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_10110,`C12T32_LLUP0_OA222X8_F_F_Z_F_10110);
		if (A && !B && C && !D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_10100,`C12T32_LLUP0_OA222X8_F_F_Z_F_10100);
		if (A && B && !C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_11010,`C12T32_LLUP0_OA222X8_F_F_Z_F_11010);
		if (!A && B && C && !D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_01100,`C12T32_LLUP0_OA222X8_F_F_Z_F_01100);
		if (!A && B && !C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_01010,`C12T32_LLUP0_OA222X8_F_F_Z_F_01010);
		if (!A && B && C && D && !E) (F +=> Z) = (`C12T32_LLUP0_OA222X8_F_R_Z_R_01110,`C12T32_LLUP0_OA222X8_F_F_Z_F_01110);


	endspecify

endmodule // C12T32_LLUP0_OA222X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA22X17_A_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X17_A_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X17_A_R_Z_R_001 0.1
`define C12T32_LLUP0_OA22X17_A_F_Z_F_001 0.1
`define C12T32_LLUP0_OA22X17_A_R_Z_R_011 0.1
`define C12T32_LLUP0_OA22X17_A_F_Z_F_011 0.1
`define C12T32_LLUP0_OA22X17_B_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X17_B_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X17_B_R_Z_R_001 0.1
`define C12T32_LLUP0_OA22X17_B_F_Z_F_001 0.1
`define C12T32_LLUP0_OA22X17_B_R_Z_R_011 0.1
`define C12T32_LLUP0_OA22X17_B_F_Z_F_011 0.1
`define C12T32_LLUP0_OA22X17_C_R_Z_R_100 0.1
`define C12T32_LLUP0_OA22X17_C_F_Z_F_100 0.1
`define C12T32_LLUP0_OA22X17_C_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X17_C_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X17_C_R_Z_R_110 0.1
`define C12T32_LLUP0_OA22X17_C_F_Z_F_110 0.1
`define C12T32_LLUP0_OA22X17_D_R_Z_R_100 0.1
`define C12T32_LLUP0_OA22X17_D_F_Z_F_100 0.1
`define C12T32_LLUP0_OA22X17_D_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X17_D_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X17_D_R_Z_R_110 0.1
`define C12T32_LLUP0_OA22X17_D_F_Z_F_110 0.1

module C12T32_LLUP0_OA22X17 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	or    U1 (INTERNAL1, A, B) ;
	or    U2 (INTERNAL2, C, D) ;
	and   #1 U3 (Z, INTERNAL1, INTERNAL2) ;



	specify

		if (!B && C && !D) (A +=> Z) = (`C12T32_LLUP0_OA22X17_A_R_Z_R_010,`C12T32_LLUP0_OA22X17_A_F_Z_F_010);
		if (!B && !C && D) (A +=> Z) = (`C12T32_LLUP0_OA22X17_A_R_Z_R_001,`C12T32_LLUP0_OA22X17_A_F_Z_F_001);
		if (!B && C && D) (A +=> Z) = (`C12T32_LLUP0_OA22X17_A_R_Z_R_011,`C12T32_LLUP0_OA22X17_A_F_Z_F_011);
		if (!A && C && !D) (B +=> Z) = (`C12T32_LLUP0_OA22X17_B_R_Z_R_010,`C12T32_LLUP0_OA22X17_B_F_Z_F_010);
		if (!A && !C && D) (B +=> Z) = (`C12T32_LLUP0_OA22X17_B_R_Z_R_001,`C12T32_LLUP0_OA22X17_B_F_Z_F_001);
		if (!A && C && D) (B +=> Z) = (`C12T32_LLUP0_OA22X17_B_R_Z_R_011,`C12T32_LLUP0_OA22X17_B_F_Z_F_011);
		if (A && !B && !D) (C +=> Z) = (`C12T32_LLUP0_OA22X17_C_R_Z_R_100,`C12T32_LLUP0_OA22X17_C_F_Z_F_100);
		if (!A && B && !D) (C +=> Z) = (`C12T32_LLUP0_OA22X17_C_R_Z_R_010,`C12T32_LLUP0_OA22X17_C_F_Z_F_010);
		if (A && B && !D) (C +=> Z) = (`C12T32_LLUP0_OA22X17_C_R_Z_R_110,`C12T32_LLUP0_OA22X17_C_F_Z_F_110);
		if (A && !B && !C) (D +=> Z) = (`C12T32_LLUP0_OA22X17_D_R_Z_R_100,`C12T32_LLUP0_OA22X17_D_F_Z_F_100);
		if (!A && B && !C) (D +=> Z) = (`C12T32_LLUP0_OA22X17_D_R_Z_R_010,`C12T32_LLUP0_OA22X17_D_F_Z_F_010);
		if (A && B && !C) (D +=> Z) = (`C12T32_LLUP0_OA22X17_D_R_Z_R_110,`C12T32_LLUP0_OA22X17_D_F_Z_F_110);


	endspecify

endmodule // C12T32_LLUP0_OA22X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OA22X8_A_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X8_A_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X8_A_R_Z_R_001 0.1
`define C12T32_LLUP0_OA22X8_A_F_Z_F_001 0.1
`define C12T32_LLUP0_OA22X8_A_R_Z_R_011 0.1
`define C12T32_LLUP0_OA22X8_A_F_Z_F_011 0.1
`define C12T32_LLUP0_OA22X8_B_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X8_B_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X8_B_R_Z_R_001 0.1
`define C12T32_LLUP0_OA22X8_B_F_Z_F_001 0.1
`define C12T32_LLUP0_OA22X8_B_R_Z_R_011 0.1
`define C12T32_LLUP0_OA22X8_B_F_Z_F_011 0.1
`define C12T32_LLUP0_OA22X8_C_R_Z_R_100 0.1
`define C12T32_LLUP0_OA22X8_C_F_Z_F_100 0.1
`define C12T32_LLUP0_OA22X8_C_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X8_C_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X8_C_R_Z_R_110 0.1
`define C12T32_LLUP0_OA22X8_C_F_Z_F_110 0.1
`define C12T32_LLUP0_OA22X8_D_R_Z_R_100 0.1
`define C12T32_LLUP0_OA22X8_D_F_Z_F_100 0.1
`define C12T32_LLUP0_OA22X8_D_R_Z_R_010 0.1
`define C12T32_LLUP0_OA22X8_D_F_Z_F_010 0.1
`define C12T32_LLUP0_OA22X8_D_R_Z_R_110 0.1
`define C12T32_LLUP0_OA22X8_D_F_Z_F_110 0.1

module C12T32_LLUP0_OA22X8 (Z, A, B, C, D);

	output Z;
	input A;
	input B;
	input C;
	input D;

	or    U1 (INTERNAL1, A, B) ;
	or    U2 (INTERNAL2, C, D) ;
	and   #1 U3 (Z, INTERNAL1, INTERNAL2) ;



	specify

		if (!B && C && !D) (A +=> Z) = (`C12T32_LLUP0_OA22X8_A_R_Z_R_010,`C12T32_LLUP0_OA22X8_A_F_Z_F_010);
		if (!B && !C && D) (A +=> Z) = (`C12T32_LLUP0_OA22X8_A_R_Z_R_001,`C12T32_LLUP0_OA22X8_A_F_Z_F_001);
		if (!B && C && D) (A +=> Z) = (`C12T32_LLUP0_OA22X8_A_R_Z_R_011,`C12T32_LLUP0_OA22X8_A_F_Z_F_011);
		if (!A && C && !D) (B +=> Z) = (`C12T32_LLUP0_OA22X8_B_R_Z_R_010,`C12T32_LLUP0_OA22X8_B_F_Z_F_010);
		if (!A && !C && D) (B +=> Z) = (`C12T32_LLUP0_OA22X8_B_R_Z_R_001,`C12T32_LLUP0_OA22X8_B_F_Z_F_001);
		if (!A && C && D) (B +=> Z) = (`C12T32_LLUP0_OA22X8_B_R_Z_R_011,`C12T32_LLUP0_OA22X8_B_F_Z_F_011);
		if (A && !B && !D) (C +=> Z) = (`C12T32_LLUP0_OA22X8_C_R_Z_R_100,`C12T32_LLUP0_OA22X8_C_F_Z_F_100);
		if (!A && B && !D) (C +=> Z) = (`C12T32_LLUP0_OA22X8_C_R_Z_R_010,`C12T32_LLUP0_OA22X8_C_F_Z_F_010);
		if (A && B && !D) (C +=> Z) = (`C12T32_LLUP0_OA22X8_C_R_Z_R_110,`C12T32_LLUP0_OA22X8_C_F_Z_F_110);
		if (A && !B && !C) (D +=> Z) = (`C12T32_LLUP0_OA22X8_D_R_Z_R_100,`C12T32_LLUP0_OA22X8_D_F_Z_F_100);
		if (!A && B && !C) (D +=> Z) = (`C12T32_LLUP0_OA22X8_D_R_Z_R_010,`C12T32_LLUP0_OA22X8_D_F_Z_F_010);
		if (A && B && !C) (D +=> Z) = (`C12T32_LLUP0_OA22X8_D_R_Z_R_110,`C12T32_LLUP0_OA22X8_D_F_Z_F_110);


	endspecify

endmodule // C12T32_LLUP0_OA22X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_OAI21X11_A_R_Z_F_01 0.1
`define C12T32_LLUP0_OAI21X11_A_F_Z_R_01 0.1
`define C12T32_LLUP0_OAI21X11_B_R_Z_F_01 0.1
`define C12T32_LLUP0_OAI21X11_B_F_Z_R_01 0.1
`define C12T32_LLUP0_OAI21X11_C_R_Z_F_01 0.1
`define C12T32_LLUP0_OAI21X11_C_F_Z_R_01 0.1
`define C12T32_LLUP0_OAI21X11_C_R_Z_F_11 0.1
`define C12T32_LLUP0_OAI21X11_C_F_Z_R_11 0.1
`define C12T32_LLUP0_OAI21X11_C_R_Z_F_10 0.1
`define C12T32_LLUP0_OAI21X11_C_F_Z_R_10 0.1

module C12T32_LLUP0_OAI21X11 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	or    U1 (INTERNAL2, A, B) ;
	and    U2 (INTERNAL1, INTERNAL2, C) ;
	not   #1 U3 (Z, INTERNAL1) ;



	specify

		if (!B && C) (A -=> Z) = (`C12T32_LLUP0_OAI21X11_A_F_Z_R_01,`C12T32_LLUP0_OAI21X11_A_R_Z_F_01);
		if (!A && C) (B -=> Z) = (`C12T32_LLUP0_OAI21X11_B_F_Z_R_01,`C12T32_LLUP0_OAI21X11_B_R_Z_F_01);
		if (!A && B) (C -=> Z) = (`C12T32_LLUP0_OAI21X11_C_F_Z_R_01,`C12T32_LLUP0_OAI21X11_C_R_Z_F_01);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_OAI21X11_C_F_Z_R_11,`C12T32_LLUP0_OAI21X11_C_R_Z_F_11);
		if (A && !B) (C -=> Z) = (`C12T32_LLUP0_OAI21X11_C_F_Z_R_10,`C12T32_LLUP0_OAI21X11_C_R_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_OAI21X11


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_PAO2X16_A_R_Z_R_01 0.1
`define C12T32_LLUP0_PAO2X16_A_F_Z_F_01 0.1
`define C12T32_LLUP0_PAO2X16_A_R_Z_R_10 0.1
`define C12T32_LLUP0_PAO2X16_A_F_Z_F_10 0.1
`define C12T32_LLUP0_PAO2X16_B_R_Z_R_01 0.1
`define C12T32_LLUP0_PAO2X16_B_F_Z_F_01 0.1
`define C12T32_LLUP0_PAO2X16_B_R_Z_R_10 0.1
`define C12T32_LLUP0_PAO2X16_B_F_Z_F_10 0.1
`define C12T32_LLUP0_PAO2X16_P_R_Z_R_01 0.1
`define C12T32_LLUP0_PAO2X16_P_F_Z_F_01 0.1
`define C12T32_LLUP0_PAO2X16_P_R_Z_R_10 0.1
`define C12T32_LLUP0_PAO2X16_P_F_Z_F_10 0.1

module C12T32_LLUP0_PAO2X16 (Z, A, B, P);

	output Z;
	input A;
	input B;
	input P;

	or    U1 (INTERNAL2, B, P) ;
	and    U2 (INTERNAL1, INTERNAL2, A) ;
	and    U3 (INTERNAL3, B, P) ;
	or   #1 U4 (Z, INTERNAL1, INTERNAL3) ;



	specify

		if (!B && P) (A +=> Z) = (`C12T32_LLUP0_PAO2X16_A_R_Z_R_01,`C12T32_LLUP0_PAO2X16_A_F_Z_F_01);
		if (B && !P) (A +=> Z) = (`C12T32_LLUP0_PAO2X16_A_R_Z_R_10,`C12T32_LLUP0_PAO2X16_A_F_Z_F_10);
		if (!A && P) (B +=> Z) = (`C12T32_LLUP0_PAO2X16_B_R_Z_R_01,`C12T32_LLUP0_PAO2X16_B_F_Z_F_01);
		if (A && !P) (B +=> Z) = (`C12T32_LLUP0_PAO2X16_B_R_Z_R_10,`C12T32_LLUP0_PAO2X16_B_F_Z_F_10);
		if (!A && B) (P +=> Z) = (`C12T32_LLUP0_PAO2X16_P_R_Z_R_01,`C12T32_LLUP0_PAO2X16_P_F_Z_F_01);
		if (A && !B) (P +=> Z) = (`C12T32_LLUP0_PAO2X16_P_R_Z_R_10,`C12T32_LLUP0_PAO2X16_P_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_PAO2X16


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_PAO2X8_A_R_Z_R_01 0.1
`define C12T32_LLUP0_PAO2X8_A_F_Z_F_01 0.1
`define C12T32_LLUP0_PAO2X8_A_R_Z_R_10 0.1
`define C12T32_LLUP0_PAO2X8_A_F_Z_F_10 0.1
`define C12T32_LLUP0_PAO2X8_B_R_Z_R_01 0.1
`define C12T32_LLUP0_PAO2X8_B_F_Z_F_01 0.1
`define C12T32_LLUP0_PAO2X8_B_R_Z_R_10 0.1
`define C12T32_LLUP0_PAO2X8_B_F_Z_F_10 0.1
`define C12T32_LLUP0_PAO2X8_P_R_Z_R_01 0.1
`define C12T32_LLUP0_PAO2X8_P_F_Z_F_01 0.1
`define C12T32_LLUP0_PAO2X8_P_R_Z_R_10 0.1
`define C12T32_LLUP0_PAO2X8_P_F_Z_F_10 0.1

module C12T32_LLUP0_PAO2X8 (Z, A, B, P);

	output Z;
	input A;
	input B;
	input P;

	or    U1 (INTERNAL2, B, P) ;
	and    U2 (INTERNAL1, INTERNAL2, A) ;
	and    U3 (INTERNAL3, B, P) ;
	or   #1 U4 (Z, INTERNAL1, INTERNAL3) ;



	specify

		if (!B && P) (A +=> Z) = (`C12T32_LLUP0_PAO2X8_A_R_Z_R_01,`C12T32_LLUP0_PAO2X8_A_F_Z_F_01);
		if (B && !P) (A +=> Z) = (`C12T32_LLUP0_PAO2X8_A_R_Z_R_10,`C12T32_LLUP0_PAO2X8_A_F_Z_F_10);
		if (!A && P) (B +=> Z) = (`C12T32_LLUP0_PAO2X8_B_R_Z_R_01,`C12T32_LLUP0_PAO2X8_B_F_Z_F_01);
		if (A && !P) (B +=> Z) = (`C12T32_LLUP0_PAO2X8_B_R_Z_R_10,`C12T32_LLUP0_PAO2X8_B_F_Z_F_10);
		if (!A && B) (P +=> Z) = (`C12T32_LLUP0_PAO2X8_P_R_Z_R_01,`C12T32_LLUP0_PAO2X8_P_F_Z_F_01);
		if (A && !B) (P +=> Z) = (`C12T32_LLUP0_PAO2X8_P_R_Z_R_10,`C12T32_LLUP0_PAO2X8_P_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_PAO2X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XNOR2X17_A_R_Z_R_1 0.1
`define C12T32_LLUP0_XNOR2X17_A_F_Z_F_1 0.1
`define C12T32_LLUP0_XNOR2X17_A_R_Z_F_0 0.1
`define C12T32_LLUP0_XNOR2X17_A_F_Z_R_0 0.1
`define C12T32_LLUP0_XNOR2X17_B_R_Z_R_1 0.1
`define C12T32_LLUP0_XNOR2X17_B_F_Z_F_1 0.1
`define C12T32_LLUP0_XNOR2X17_B_R_Z_F_0 0.1
`define C12T32_LLUP0_XNOR2X17_B_F_Z_R_0 0.1

module C12T32_LLUP0_XNOR2X17 (Z, A, B);

	output Z;
	input A;
	input B;

	xor    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A +=> Z) = (`C12T32_LLUP0_XNOR2X17_A_R_Z_R_1,`C12T32_LLUP0_XNOR2X17_A_F_Z_F_1);
		if (!B) (A -=> Z) = (`C12T32_LLUP0_XNOR2X17_A_F_Z_R_0,`C12T32_LLUP0_XNOR2X17_A_R_Z_F_0);
		if (A) (B +=> Z) = (`C12T32_LLUP0_XNOR2X17_B_R_Z_R_1,`C12T32_LLUP0_XNOR2X17_B_F_Z_F_1);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_XNOR2X17_B_F_Z_R_0,`C12T32_LLUP0_XNOR2X17_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_XNOR2X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XNOR2X8_A_R_Z_R_1 0.1
`define C12T32_LLUP0_XNOR2X8_A_F_Z_F_1 0.1
`define C12T32_LLUP0_XNOR2X8_A_R_Z_F_0 0.1
`define C12T32_LLUP0_XNOR2X8_A_F_Z_R_0 0.1
`define C12T32_LLUP0_XNOR2X8_B_R_Z_R_1 0.1
`define C12T32_LLUP0_XNOR2X8_B_F_Z_F_1 0.1
`define C12T32_LLUP0_XNOR2X8_B_R_Z_F_0 0.1
`define C12T32_LLUP0_XNOR2X8_B_F_Z_R_0 0.1

module C12T32_LLUP0_XNOR2X8 (Z, A, B);

	output Z;
	input A;
	input B;

	xor    U1 (INTERNAL1, A, B) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B) (A +=> Z) = (`C12T32_LLUP0_XNOR2X8_A_R_Z_R_1,`C12T32_LLUP0_XNOR2X8_A_F_Z_F_1);
		if (!B) (A -=> Z) = (`C12T32_LLUP0_XNOR2X8_A_F_Z_R_0,`C12T32_LLUP0_XNOR2X8_A_R_Z_F_0);
		if (A) (B +=> Z) = (`C12T32_LLUP0_XNOR2X8_B_R_Z_R_1,`C12T32_LLUP0_XNOR2X8_B_F_Z_F_1);
		if (!A) (B -=> Z) = (`C12T32_LLUP0_XNOR2X8_B_F_Z_R_0,`C12T32_LLUP0_XNOR2X8_B_R_Z_F_0);


	endspecify

endmodule // C12T32_LLUP0_XNOR2X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XNOR3X16_A_R_Z_F_11 0.1
`define C12T32_LLUP0_XNOR3X16_A_F_Z_R_11 0.1
`define C12T32_LLUP0_XNOR3X16_A_R_Z_F_00 0.1
`define C12T32_LLUP0_XNOR3X16_A_F_Z_R_00 0.1
`define C12T32_LLUP0_XNOR3X16_A_R_Z_R_01 0.1
`define C12T32_LLUP0_XNOR3X16_A_F_Z_F_01 0.1
`define C12T32_LLUP0_XNOR3X16_A_R_Z_R_10 0.1
`define C12T32_LLUP0_XNOR3X16_A_F_Z_F_10 0.1
`define C12T32_LLUP0_XNOR3X16_B_R_Z_F_11 0.1
`define C12T32_LLUP0_XNOR3X16_B_F_Z_R_11 0.1
`define C12T32_LLUP0_XNOR3X16_B_R_Z_F_00 0.1
`define C12T32_LLUP0_XNOR3X16_B_F_Z_R_00 0.1
`define C12T32_LLUP0_XNOR3X16_B_R_Z_R_01 0.1
`define C12T32_LLUP0_XNOR3X16_B_F_Z_F_01 0.1
`define C12T32_LLUP0_XNOR3X16_B_R_Z_R_10 0.1
`define C12T32_LLUP0_XNOR3X16_B_F_Z_F_10 0.1
`define C12T32_LLUP0_XNOR3X16_C_R_Z_F_11 0.1
`define C12T32_LLUP0_XNOR3X16_C_F_Z_R_11 0.1
`define C12T32_LLUP0_XNOR3X16_C_R_Z_F_00 0.1
`define C12T32_LLUP0_XNOR3X16_C_F_Z_R_00 0.1
`define C12T32_LLUP0_XNOR3X16_C_R_Z_R_01 0.1
`define C12T32_LLUP0_XNOR3X16_C_F_Z_F_01 0.1
`define C12T32_LLUP0_XNOR3X16_C_R_Z_R_10 0.1
`define C12T32_LLUP0_XNOR3X16_C_F_Z_F_10 0.1

module C12T32_LLUP0_XNOR3X16 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	xor    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_XNOR3X16_A_F_Z_R_11,`C12T32_LLUP0_XNOR3X16_A_R_Z_F_11);
		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_XNOR3X16_A_F_Z_R_00,`C12T32_LLUP0_XNOR3X16_A_R_Z_F_00);
		if (!B && C) (A +=> Z) = (`C12T32_LLUP0_XNOR3X16_A_R_Z_R_01,`C12T32_LLUP0_XNOR3X16_A_F_Z_F_01);
		if (B && !C) (A +=> Z) = (`C12T32_LLUP0_XNOR3X16_A_R_Z_R_10,`C12T32_LLUP0_XNOR3X16_A_F_Z_F_10);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_XNOR3X16_B_F_Z_R_11,`C12T32_LLUP0_XNOR3X16_B_R_Z_F_11);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_XNOR3X16_B_F_Z_R_00,`C12T32_LLUP0_XNOR3X16_B_R_Z_F_00);
		if (!A && C) (B +=> Z) = (`C12T32_LLUP0_XNOR3X16_B_R_Z_R_01,`C12T32_LLUP0_XNOR3X16_B_F_Z_F_01);
		if (A && !C) (B +=> Z) = (`C12T32_LLUP0_XNOR3X16_B_R_Z_R_10,`C12T32_LLUP0_XNOR3X16_B_F_Z_F_10);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_XNOR3X16_C_F_Z_R_11,`C12T32_LLUP0_XNOR3X16_C_R_Z_F_11);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_XNOR3X16_C_F_Z_R_00,`C12T32_LLUP0_XNOR3X16_C_R_Z_F_00);
		if (!A && B) (C +=> Z) = (`C12T32_LLUP0_XNOR3X16_C_R_Z_R_01,`C12T32_LLUP0_XNOR3X16_C_F_Z_F_01);
		if (A && !B) (C +=> Z) = (`C12T32_LLUP0_XNOR3X16_C_R_Z_R_10,`C12T32_LLUP0_XNOR3X16_C_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_XNOR3X16


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XNOR3X8_A_R_Z_F_11 0.1
`define C12T32_LLUP0_XNOR3X8_A_F_Z_R_11 0.1
`define C12T32_LLUP0_XNOR3X8_A_R_Z_F_00 0.1
`define C12T32_LLUP0_XNOR3X8_A_F_Z_R_00 0.1
`define C12T32_LLUP0_XNOR3X8_A_R_Z_R_01 0.1
`define C12T32_LLUP0_XNOR3X8_A_F_Z_F_01 0.1
`define C12T32_LLUP0_XNOR3X8_A_R_Z_R_10 0.1
`define C12T32_LLUP0_XNOR3X8_A_F_Z_F_10 0.1
`define C12T32_LLUP0_XNOR3X8_B_R_Z_F_11 0.1
`define C12T32_LLUP0_XNOR3X8_B_F_Z_R_11 0.1
`define C12T32_LLUP0_XNOR3X8_B_R_Z_F_00 0.1
`define C12T32_LLUP0_XNOR3X8_B_F_Z_R_00 0.1
`define C12T32_LLUP0_XNOR3X8_B_R_Z_R_01 0.1
`define C12T32_LLUP0_XNOR3X8_B_F_Z_F_01 0.1
`define C12T32_LLUP0_XNOR3X8_B_R_Z_R_10 0.1
`define C12T32_LLUP0_XNOR3X8_B_F_Z_F_10 0.1
`define C12T32_LLUP0_XNOR3X8_C_R_Z_F_11 0.1
`define C12T32_LLUP0_XNOR3X8_C_F_Z_R_11 0.1
`define C12T32_LLUP0_XNOR3X8_C_R_Z_F_00 0.1
`define C12T32_LLUP0_XNOR3X8_C_F_Z_R_00 0.1
`define C12T32_LLUP0_XNOR3X8_C_R_Z_R_01 0.1
`define C12T32_LLUP0_XNOR3X8_C_F_Z_F_01 0.1
`define C12T32_LLUP0_XNOR3X8_C_R_Z_R_10 0.1
`define C12T32_LLUP0_XNOR3X8_C_F_Z_F_10 0.1

module C12T32_LLUP0_XNOR3X8 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	xor    U1 (INTERNAL1, A, B, C) ;
	not   #1 U2 (Z, INTERNAL1) ;



	specify

		if (B && C) (A -=> Z) = (`C12T32_LLUP0_XNOR3X8_A_F_Z_R_11,`C12T32_LLUP0_XNOR3X8_A_R_Z_F_11);
		if (!B && !C) (A -=> Z) = (`C12T32_LLUP0_XNOR3X8_A_F_Z_R_00,`C12T32_LLUP0_XNOR3X8_A_R_Z_F_00);
		if (!B && C) (A +=> Z) = (`C12T32_LLUP0_XNOR3X8_A_R_Z_R_01,`C12T32_LLUP0_XNOR3X8_A_F_Z_F_01);
		if (B && !C) (A +=> Z) = (`C12T32_LLUP0_XNOR3X8_A_R_Z_R_10,`C12T32_LLUP0_XNOR3X8_A_F_Z_F_10);
		if (A && C) (B -=> Z) = (`C12T32_LLUP0_XNOR3X8_B_F_Z_R_11,`C12T32_LLUP0_XNOR3X8_B_R_Z_F_11);
		if (!A && !C) (B -=> Z) = (`C12T32_LLUP0_XNOR3X8_B_F_Z_R_00,`C12T32_LLUP0_XNOR3X8_B_R_Z_F_00);
		if (!A && C) (B +=> Z) = (`C12T32_LLUP0_XNOR3X8_B_R_Z_R_01,`C12T32_LLUP0_XNOR3X8_B_F_Z_F_01);
		if (A && !C) (B +=> Z) = (`C12T32_LLUP0_XNOR3X8_B_R_Z_R_10,`C12T32_LLUP0_XNOR3X8_B_F_Z_F_10);
		if (A && B) (C -=> Z) = (`C12T32_LLUP0_XNOR3X8_C_F_Z_R_11,`C12T32_LLUP0_XNOR3X8_C_R_Z_F_11);
		if (!A && !B) (C -=> Z) = (`C12T32_LLUP0_XNOR3X8_C_F_Z_R_00,`C12T32_LLUP0_XNOR3X8_C_R_Z_F_00);
		if (!A && B) (C +=> Z) = (`C12T32_LLUP0_XNOR3X8_C_R_Z_R_01,`C12T32_LLUP0_XNOR3X8_C_F_Z_F_01);
		if (A && !B) (C +=> Z) = (`C12T32_LLUP0_XNOR3X8_C_R_Z_R_10,`C12T32_LLUP0_XNOR3X8_C_F_Z_F_10);


	endspecify

endmodule // C12T32_LLUP0_XNOR3X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XOR2X16_A_R_Z_R_0 0.1
`define C12T32_LLUP0_XOR2X16_A_F_Z_F_0 0.1
`define C12T32_LLUP0_XOR2X16_A_R_Z_F_1 0.1
`define C12T32_LLUP0_XOR2X16_A_F_Z_R_1 0.1
`define C12T32_LLUP0_XOR2X16_B_R_Z_R_0 0.1
`define C12T32_LLUP0_XOR2X16_B_F_Z_F_0 0.1
`define C12T32_LLUP0_XOR2X16_B_R_Z_F_1 0.1
`define C12T32_LLUP0_XOR2X16_B_F_Z_R_1 0.1

module C12T32_LLUP0_XOR2X16 (Z, A, B);

	output Z;
	input A;
	input B;

	xor   #1 U1 (Z, A, B) ;



	specify

		if (!B) (A +=> Z) = (`C12T32_LLUP0_XOR2X16_A_R_Z_R_0,`C12T32_LLUP0_XOR2X16_A_F_Z_F_0);
		if (B) (A -=> Z) = (`C12T32_LLUP0_XOR2X16_A_F_Z_R_1,`C12T32_LLUP0_XOR2X16_A_R_Z_F_1);
		if (!A) (B +=> Z) = (`C12T32_LLUP0_XOR2X16_B_R_Z_R_0,`C12T32_LLUP0_XOR2X16_B_F_Z_F_0);
		if (A) (B -=> Z) = (`C12T32_LLUP0_XOR2X16_B_F_Z_R_1,`C12T32_LLUP0_XOR2X16_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_XOR2X16


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XOR2X4_A_R_Z_R_0 0.1
`define C12T32_LLUP0_XOR2X4_A_F_Z_F_0 0.1
`define C12T32_LLUP0_XOR2X4_A_R_Z_F_1 0.1
`define C12T32_LLUP0_XOR2X4_A_F_Z_R_1 0.1
`define C12T32_LLUP0_XOR2X4_B_R_Z_R_0 0.1
`define C12T32_LLUP0_XOR2X4_B_F_Z_F_0 0.1
`define C12T32_LLUP0_XOR2X4_B_R_Z_F_1 0.1
`define C12T32_LLUP0_XOR2X4_B_F_Z_R_1 0.1

module C12T32_LLUP0_XOR2X4 (Z, A, B);

	output Z;
	input A;
	input B;

	xor   #1 U1 (Z, A, B) ;



	specify

		if (!B) (A +=> Z) = (`C12T32_LLUP0_XOR2X4_A_R_Z_R_0,`C12T32_LLUP0_XOR2X4_A_F_Z_F_0);
		if (B) (A -=> Z) = (`C12T32_LLUP0_XOR2X4_A_F_Z_R_1,`C12T32_LLUP0_XOR2X4_A_R_Z_F_1);
		if (!A) (B +=> Z) = (`C12T32_LLUP0_XOR2X4_B_R_Z_R_0,`C12T32_LLUP0_XOR2X4_B_F_Z_F_0);
		if (A) (B -=> Z) = (`C12T32_LLUP0_XOR2X4_B_F_Z_R_1,`C12T32_LLUP0_XOR2X4_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_XOR2X4


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XOR2X8_A_R_Z_R_0 0.1
`define C12T32_LLUP0_XOR2X8_A_F_Z_F_0 0.1
`define C12T32_LLUP0_XOR2X8_A_R_Z_F_1 0.1
`define C12T32_LLUP0_XOR2X8_A_F_Z_R_1 0.1
`define C12T32_LLUP0_XOR2X8_B_R_Z_R_0 0.1
`define C12T32_LLUP0_XOR2X8_B_F_Z_F_0 0.1
`define C12T32_LLUP0_XOR2X8_B_R_Z_F_1 0.1
`define C12T32_LLUP0_XOR2X8_B_F_Z_R_1 0.1

module C12T32_LLUP0_XOR2X8 (Z, A, B);

	output Z;
	input A;
	input B;

	xor   #1 U1 (Z, A, B) ;



	specify

		if (!B) (A +=> Z) = (`C12T32_LLUP0_XOR2X8_A_R_Z_R_0,`C12T32_LLUP0_XOR2X8_A_F_Z_F_0);
		if (B) (A -=> Z) = (`C12T32_LLUP0_XOR2X8_A_F_Z_R_1,`C12T32_LLUP0_XOR2X8_A_R_Z_F_1);
		if (!A) (B +=> Z) = (`C12T32_LLUP0_XOR2X8_B_R_Z_R_0,`C12T32_LLUP0_XOR2X8_B_F_Z_F_0);
		if (A) (B -=> Z) = (`C12T32_LLUP0_XOR2X8_B_F_Z_R_1,`C12T32_LLUP0_XOR2X8_B_R_Z_F_1);


	endspecify

endmodule // C12T32_LLUP0_XOR2X8


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XOR3X17_A_R_Z_F_10 0.1
`define C12T32_LLUP0_XOR3X17_A_F_Z_R_10 0.1
`define C12T32_LLUP0_XOR3X17_A_R_Z_F_01 0.1
`define C12T32_LLUP0_XOR3X17_A_F_Z_R_01 0.1
`define C12T32_LLUP0_XOR3X17_A_R_Z_R_00 0.1
`define C12T32_LLUP0_XOR3X17_A_F_Z_F_00 0.1
`define C12T32_LLUP0_XOR3X17_A_R_Z_R_11 0.1
`define C12T32_LLUP0_XOR3X17_A_F_Z_F_11 0.1
`define C12T32_LLUP0_XOR3X17_B_R_Z_F_10 0.1
`define C12T32_LLUP0_XOR3X17_B_F_Z_R_10 0.1
`define C12T32_LLUP0_XOR3X17_B_R_Z_F_01 0.1
`define C12T32_LLUP0_XOR3X17_B_F_Z_R_01 0.1
`define C12T32_LLUP0_XOR3X17_B_R_Z_R_00 0.1
`define C12T32_LLUP0_XOR3X17_B_F_Z_F_00 0.1
`define C12T32_LLUP0_XOR3X17_B_R_Z_R_11 0.1
`define C12T32_LLUP0_XOR3X17_B_F_Z_F_11 0.1
`define C12T32_LLUP0_XOR3X17_C_R_Z_F_10 0.1
`define C12T32_LLUP0_XOR3X17_C_F_Z_R_10 0.1
`define C12T32_LLUP0_XOR3X17_C_R_Z_F_01 0.1
`define C12T32_LLUP0_XOR3X17_C_F_Z_R_01 0.1
`define C12T32_LLUP0_XOR3X17_C_R_Z_R_00 0.1
`define C12T32_LLUP0_XOR3X17_C_F_Z_F_00 0.1
`define C12T32_LLUP0_XOR3X17_C_R_Z_R_11 0.1
`define C12T32_LLUP0_XOR3X17_C_F_Z_F_11 0.1

module C12T32_LLUP0_XOR3X17 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	xor   #1 U1 (Z, A, B, C) ;



	specify

		if (B && !C) (A -=> Z) = (`C12T32_LLUP0_XOR3X17_A_F_Z_R_10,`C12T32_LLUP0_XOR3X17_A_R_Z_F_10);
		if (!B && C) (A -=> Z) = (`C12T32_LLUP0_XOR3X17_A_F_Z_R_01,`C12T32_LLUP0_XOR3X17_A_R_Z_F_01);
		if (!B && !C) (A +=> Z) = (`C12T32_LLUP0_XOR3X17_A_R_Z_R_00,`C12T32_LLUP0_XOR3X17_A_F_Z_F_00);
		if (B && C) (A +=> Z) = (`C12T32_LLUP0_XOR3X17_A_R_Z_R_11,`C12T32_LLUP0_XOR3X17_A_F_Z_F_11);
		if (A && !C) (B -=> Z) = (`C12T32_LLUP0_XOR3X17_B_F_Z_R_10,`C12T32_LLUP0_XOR3X17_B_R_Z_F_10);
		if (!A && C) (B -=> Z) = (`C12T32_LLUP0_XOR3X17_B_F_Z_R_01,`C12T32_LLUP0_XOR3X17_B_R_Z_F_01);
		if (!A && !C) (B +=> Z) = (`C12T32_LLUP0_XOR3X17_B_R_Z_R_00,`C12T32_LLUP0_XOR3X17_B_F_Z_F_00);
		if (A && C) (B +=> Z) = (`C12T32_LLUP0_XOR3X17_B_R_Z_R_11,`C12T32_LLUP0_XOR3X17_B_F_Z_F_11);
		if (A && !B) (C -=> Z) = (`C12T32_LLUP0_XOR3X17_C_F_Z_R_10,`C12T32_LLUP0_XOR3X17_C_R_Z_F_10);
		if (!A && B) (C -=> Z) = (`C12T32_LLUP0_XOR3X17_C_F_Z_R_01,`C12T32_LLUP0_XOR3X17_C_R_Z_F_01);
		if (!A && !B) (C +=> Z) = (`C12T32_LLUP0_XOR3X17_C_R_Z_R_00,`C12T32_LLUP0_XOR3X17_C_F_Z_F_00);
		if (A && B) (C +=> Z) = (`C12T32_LLUP0_XOR3X17_C_R_Z_R_11,`C12T32_LLUP0_XOR3X17_C_F_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_XOR3X17


`endcelldefine
`celldefine
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 1ps
   `delay_mode_path
`endif

`define C12T32_LLUP0_XOR3X8_A_R_Z_F_10 0.1
`define C12T32_LLUP0_XOR3X8_A_F_Z_R_10 0.1
`define C12T32_LLUP0_XOR3X8_A_R_Z_F_01 0.1
`define C12T32_LLUP0_XOR3X8_A_F_Z_R_01 0.1
`define C12T32_LLUP0_XOR3X8_A_R_Z_R_00 0.1
`define C12T32_LLUP0_XOR3X8_A_F_Z_F_00 0.1
`define C12T32_LLUP0_XOR3X8_A_R_Z_R_11 0.1
`define C12T32_LLUP0_XOR3X8_A_F_Z_F_11 0.1
`define C12T32_LLUP0_XOR3X8_B_R_Z_F_10 0.1
`define C12T32_LLUP0_XOR3X8_B_F_Z_R_10 0.1
`define C12T32_LLUP0_XOR3X8_B_R_Z_F_01 0.1
`define C12T32_LLUP0_XOR3X8_B_F_Z_R_01 0.1
`define C12T32_LLUP0_XOR3X8_B_R_Z_R_00 0.1
`define C12T32_LLUP0_XOR3X8_B_F_Z_F_00 0.1
`define C12T32_LLUP0_XOR3X8_B_R_Z_R_11 0.1
`define C12T32_LLUP0_XOR3X8_B_F_Z_F_11 0.1
`define C12T32_LLUP0_XOR3X8_C_R_Z_F_10 0.1
`define C12T32_LLUP0_XOR3X8_C_F_Z_R_10 0.1
`define C12T32_LLUP0_XOR3X8_C_R_Z_F_01 0.1
`define C12T32_LLUP0_XOR3X8_C_F_Z_R_01 0.1
`define C12T32_LLUP0_XOR3X8_C_R_Z_R_00 0.1
`define C12T32_LLUP0_XOR3X8_C_F_Z_F_00 0.1
`define C12T32_LLUP0_XOR3X8_C_R_Z_R_11 0.1
`define C12T32_LLUP0_XOR3X8_C_F_Z_F_11 0.1

module C12T32_LLUP0_XOR3X8 (Z, A, B, C);

	output Z;
	input A;
	input B;
	input C;

	xor   #1 U1 (Z, A, B, C) ;



	specify

		if (B && !C) (A -=> Z) = (`C12T32_LLUP0_XOR3X8_A_F_Z_R_10,`C12T32_LLUP0_XOR3X8_A_R_Z_F_10);
		if (!B && C) (A -=> Z) = (`C12T32_LLUP0_XOR3X8_A_F_Z_R_01,`C12T32_LLUP0_XOR3X8_A_R_Z_F_01);
		if (!B && !C) (A +=> Z) = (`C12T32_LLUP0_XOR3X8_A_R_Z_R_00,`C12T32_LLUP0_XOR3X8_A_F_Z_F_00);
		if (B && C) (A +=> Z) = (`C12T32_LLUP0_XOR3X8_A_R_Z_R_11,`C12T32_LLUP0_XOR3X8_A_F_Z_F_11);
		if (A && !C) (B -=> Z) = (`C12T32_LLUP0_XOR3X8_B_F_Z_R_10,`C12T32_LLUP0_XOR3X8_B_R_Z_F_10);
		if (!A && C) (B -=> Z) = (`C12T32_LLUP0_XOR3X8_B_F_Z_R_01,`C12T32_LLUP0_XOR3X8_B_R_Z_F_01);
		if (!A && !C) (B +=> Z) = (`C12T32_LLUP0_XOR3X8_B_R_Z_R_00,`C12T32_LLUP0_XOR3X8_B_F_Z_F_00);
		if (A && C) (B +=> Z) = (`C12T32_LLUP0_XOR3X8_B_R_Z_R_11,`C12T32_LLUP0_XOR3X8_B_F_Z_F_11);
		if (A && !B) (C -=> Z) = (`C12T32_LLUP0_XOR3X8_C_F_Z_R_10,`C12T32_LLUP0_XOR3X8_C_R_Z_F_10);
		if (!A && B) (C -=> Z) = (`C12T32_LLUP0_XOR3X8_C_F_Z_R_01,`C12T32_LLUP0_XOR3X8_C_R_Z_F_01);
		if (!A && !B) (C +=> Z) = (`C12T32_LLUP0_XOR3X8_C_R_Z_R_00,`C12T32_LLUP0_XOR3X8_C_F_Z_F_00);
		if (A && B) (C +=> Z) = (`C12T32_LLUP0_XOR3X8_C_R_Z_R_11,`C12T32_LLUP0_XOR3X8_C_F_Z_F_11);


	endspecify

endmodule // C12T32_LLUP0_XOR3X8


`endcelldefine

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive
primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive

primitive U_POWER (Z, Z_NOPWR, GND_FINAL, VDD_FINAL);
        output Z;
        input  Z_NOPWR, GND_FINAL, VDD_FINAL;

        table
        //Z_NOPWR       GND_FINAL       VDD_FINAL        : Z
         0      1       1 :      0 ;
         1      1       1 :      1 ;
         X      1       1 :      X ;

        endtable

endprimitive


