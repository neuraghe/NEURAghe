`include "pulp_interfaces.sv"

module noc_interconnect_wrap
#(
   parameter AXI_ADDR_WIDTH = 32,
   parameter AXI_DATA_WIDTH = 64,
   parameter AXI_ID_WIDTH   = 4,
   parameter AXI_USER_WIDTH = 6
)
(
    input  logic                clk,
    input  logic                rst,

    AXI_BUS.Master              data_master_CL0,
    AXI_BUS.Master              instr_master_CL0,
    AXI_BUS.Slave               data_slave_CL0,

    AXI_BUS.Master              data_master_CL1,
    AXI_BUS.Master              instr_master_CL1,
    AXI_BUS.Slave               data_slave_CL1,

    AXI_BUS.Master              data_master_CL2,
    AXI_BUS.Master              instr_master_CL2,
    AXI_BUS.Slave               data_slave_CL2,

    AXI_BUS.Master              data_master_CL3,
    AXI_BUS.Master              instr_master_CL3,
    AXI_BUS.Slave               data_slave_CL3,

    AXI_BUS.Master              data_master_L2_MEM,
    AXI_BUS.Slave               data_slave_EXT
);





noc_interconnect noc_interconnect_i
(
     .clk                 ( clk                       ), 
     .rst                 ( rst                       ), 

     .AWID_in_MD_CL0      ( data_master_CL0.aw_id     ),
     .AWADDR_in_MD_CL0    ( data_master_CL0.aw_addr   ),
     .AWLEN_in_MD_CL0     ( data_master_CL0.aw_len    ),
     .AWSIZE_in_MD_CL0    ( data_master_CL0.aw_size   ),
     .AWBURST_in_MD_CL0   ( data_master_CL0.aw_burst  ),
     .AWLOCK_in_MD_CL0    ( {1'b0, data_master_CL0.aw_lock}   ),
     .AWCACHE_in_MD_CL0   ( data_master_CL0.aw_cache  ),
     .AWPROT_in_MD_CL0    ( data_master_CL0.aw_prot   ),
     .AWVALID_in_MD_CL0   ( data_master_CL0.aw_valid  ),
     .AWREADY_out_MD_CL0  ( data_master_CL0.aw_ready  ),
     .WID_in_MD_CL0       ( '0                        ),
     .WDATA_in_MD_CL0     ( data_master_CL0.w_data    ),
     .WSTRB_in_MD_CL0     ( data_master_CL0.w_strb    ),
     .WLAST_in_MD_CL0     ( data_master_CL0.w_last    ),
     .WVALID_in_MD_CL0    ( data_master_CL0.w_valid   ),
     .WREADY_out_MD_CL0   ( data_master_CL0.w_ready   ),
     
     .ARID_in_MD_CL0      ( data_master_CL0.ar_id     ),
     .ARADDR_in_MD_CL0    ( data_master_CL0.ar_addr   ),
     .ARLEN_in_MD_CL0     ( data_master_CL0.ar_len    ),
     .ARSIZE_in_MD_CL0    ( data_master_CL0.ar_size   ),
     .ARBURST_in_MD_CL0   ( data_master_CL0.ar_burst  ),
     .ARLOCK_in_MD_CL0    ( {1'b0, data_master_CL0.ar_lock }  ),
     .ARCACHE_in_MD_CL0   ( data_master_CL0.ar_cache  ),
     .ARPROT_in_MD_CL0    ( data_master_CL0.ar_prot   ),
     .ARVALID_in_MD_CL0   ( data_master_CL0.ar_valid  ),
     .ARREADY_out_MD_CL0  ( data_master_CL0.ar_ready  ),

     .RID_out_MD_CL0      ( data_master_CL0.r_id      ),
     .RDATA_out_MD_CL0    ( data_master_CL0.r_data    ),
     .RRESP_out_MD_CL0    ( data_master_CL0.r_resp    ),
     .RLAST_out_MD_CL0    ( data_master_CL0.r_last    ),
     .RVALID_out_MD_CL0   ( data_master_CL0.r_valid   ),
     .RREADY_in_MD_CL0    ( data_master_CL0.r_ready   ),
     .BID_out_MD_CL0      ( data_master_CL0.b_id      ),
     .BRESP_out_MD_CL0    ( data_master_CL0.b_resp    ),
     .BVALID_out_MD_CL0   ( data_master_CL0.b_valid   ),
     .BREADY_in_MD_CL0    ( data_master_CL0.b_ready   ),
     .init_div_MD_CL0     ( 1                         ),

     .AWID_out_SD_CL0      ( data_slave_CL0.aw_id    ),
     .AWADDR_out_SD_CL0    ( data_slave_CL0.aw_addr  ),
     .AWLEN_out_SD_CL0     ( data_slave_CL0.aw_len   ),
     .AWSIZE_out_SD_CL0    ( data_slave_CL0.aw_size  ),
     .AWBURST_out_SD_CL0   ( data_slave_CL0.aw_burst ),
     .AWLOCK_out_SD_CL0    ( {tmp0,data_slave_CL0.aw_lock}  ),
     .AWCACHE_out_SD_CL0   ( data_slave_CL0.aw_cache ),
     .AWPROT_out_SD_CL0    ( data_slave_CL0.aw_prot  ),
     .AWVALID_out_SD_CL0   ( data_slave_CL0.aw_valid ),
     .AWREADY_in_SD_CL0    ( data_slave_CL0.aw_ready ),
     .WID_out_SD_CL0       (                         ),
     .WDATA_out_SD_CL0     ( data_slave_CL0.w_data   ),
     .WSTRB_out_SD_CL0     ( data_slave_CL0.w_strb   ),
     .WLAST_out_SD_CL0     ( data_slave_CL0.w_last   ),
     .WVALID_out_SD_CL0    ( data_slave_CL0.w_valid  ),
     .WREADY_in_SD_CL0     ( data_slave_CL0.w_ready  ),
     .ARID_out_SD_CL0      ( data_slave_CL0.ar_id    ),
     .ARADDR_out_SD_CL0    ( data_slave_CL0.ar_addr  ),
     .ARLEN_out_SD_CL0     ( data_slave_CL0.ar_len   ),
     .ARSIZE_out_SD_CL0    ( data_slave_CL0.ar_size  ),
     .ARBURST_out_SD_CL0   ( data_slave_CL0.ar_burst ),
     .ARLOCK_out_SD_CL0    ( {tmp1, data_slave_CL0.ar_lock}  ),
     .ARCACHE_out_SD_CL0   ( data_slave_CL0.ar_cache ),
     .ARPROT_out_SD_CL0    ( data_slave_CL0.ar_prot  ),
     .ARVALID_out_SD_CL0   ( data_slave_CL0.ar_valid ),
     .ARREADY_in_SD_CL0    ( data_slave_CL0.ar_ready ),
     .RID_in_SD_CL0        ( data_slave_CL0.r_id     ),
     .RDATA_in_SD_CL0      ( data_slave_CL0.r_data   ),
     .RRESP_in_SD_CL0      ( data_slave_CL0.r_resp   ),
     .RLAST_in_SD_CL0      ( data_slave_CL0.r_last   ),
     .RVALID_in_SD_CL0     ( data_slave_CL0.r_valid  ),
     .RREADY_out_SD_CL0    ( data_slave_CL0.r_ready  ),
     .BID_in_SD_CL0        ( data_slave_CL0.b_id     ),
     .BRESP_in_SD_CL0      ( data_slave_CL0.b_resp   ),
     .BVALID_in_SD_CL0     ( data_slave_CL0.b_valid  ),
     .BREADY_out_SD_CL0    ( data_slave_CL0.b_ready  ),
     .target_div_SD_CL0    ( 1                       ),

     .AWID_in_MI_CL0       ( instr_master_CL0.aw_id    ),
     .AWADDR_in_MI_CL0     ( instr_master_CL0.aw_addr  ),
     .AWLEN_in_MI_CL0      ( instr_master_CL0.aw_len   ),
     .AWSIZE_in_MI_CL0     ( instr_master_CL0.aw_size  ),
     .AWBURST_in_MI_CL0    ( instr_master_CL0.aw_burst ),
     .AWLOCK_in_MI_CL0     ( {1'b0, instr_master_CL0.aw_lock } ),
     .AWCACHE_in_MI_CL0    ( instr_master_CL0.aw_cache ),
     .AWPROT_in_MI_CL0     ( instr_master_CL0.aw_prot  ),
     .AWVALID_in_MI_CL0    ( instr_master_CL0.aw_valid ),
     .AWREADY_out_MI_CL0   ( instr_master_CL0.aw_ready ),
     .WID_in_MI_CL0        (                           ),
     .WDATA_in_MI_CL0      ( instr_master_CL0.w_data   ),
     .WSTRB_in_MI_CL0      ( instr_master_CL0.w_strb   ),
     .WLAST_in_MI_CL0      ( instr_master_CL0.w_last   ),
     .WVALID_in_MI_CL0     ( instr_master_CL0.w_valid  ),
     .WREADY_out_MI_CL0    ( instr_master_CL0.w_ready  ),
     .ARID_in_MI_CL0       ( instr_master_CL0.ar_id    ),
     .ARADDR_in_MI_CL0     ( instr_master_CL0.ar_addr  ),
     .ARLEN_in_MI_CL0      ( instr_master_CL0.ar_len   ),
     .ARSIZE_in_MI_CL0     ( instr_master_CL0.ar_size  ),
     .ARBURST_in_MI_CL0    ( instr_master_CL0.ar_burst ),
     .ARLOCK_in_MI_CL0     ( {1'b0, instr_master_CL0.ar_lock } ),
     .ARCACHE_in_MI_CL0    ( instr_master_CL0.ar_cache ),
     .ARPROT_in_MI_CL0     ( instr_master_CL0.ar_prot  ),
     .ARVALID_in_MI_CL0    ( instr_master_CL0.ar_valid ),
     .ARREADY_out_MI_CL0   ( instr_master_CL0.ar_ready ),
     .RID_out_MI_CL0       ( instr_master_CL0.r_id     ),
     .RDATA_out_MI_CL0     ( instr_master_CL0.r_data   ),
     .RRESP_out_MI_CL0     ( instr_master_CL0.r_resp   ),
     .RLAST_out_MI_CL0     ( instr_master_CL0.r_last   ),
     .RVALID_out_MI_CL0    ( instr_master_CL0.r_valid  ),
     .RREADY_in_MI_CL0     ( instr_master_CL0.r_ready  ),
     .BID_out_MI_CL0       ( instr_master_CL0.b_id     ),
     .BRESP_out_MI_CL0     ( instr_master_CL0.b_resp   ),
     .BVALID_out_MI_CL0    ( instr_master_CL0.b_valid  ),
     .BREADY_in_MI_CL0     ( instr_master_CL0.b_ready  ),
     .init_div_MI_CL0      ( 1                        ),

     .AWID_in_MD_CL1       ( data_master_CL1.aw_id    ),
     .AWADDR_in_MD_CL1     ( data_master_CL1.aw_addr  ),
     .AWLEN_in_MD_CL1      ( data_master_CL1.aw_len   ),
     .AWSIZE_in_MD_CL1     ( data_master_CL1.aw_size  ),
     .AWBURST_in_MD_CL1    ( data_master_CL1.aw_burst ),
     .AWLOCK_in_MD_CL1     ( data_master_CL1.aw_lock  ),
     .AWCACHE_in_MD_CL1    ( data_master_CL1.aw_cache ),
     .AWPROT_in_MD_CL1     ( data_master_CL1.aw_prot  ),
     .AWVALID_in_MD_CL1    ( data_master_CL1.aw_valid ),
     .AWREADY_out_MD_CL1   ( data_master_CL1.aw_ready ),
     .WID_in_MD_CL1        ( '0                       ),
     .WDATA_in_MD_CL1      ( data_master_CL1.w_data   ),
     .WSTRB_in_MD_CL1      ( data_master_CL1.w_strb   ),
     .WLAST_in_MD_CL1      ( data_master_CL1.w_last   ),
     .WVALID_in_MD_CL1     ( data_master_CL1.w_valid  ),
     .WREADY_out_MD_CL1    ( data_master_CL1.w_ready  ),
     .ARID_in_MD_CL1       ( data_master_CL1.ar_id    ),
     .ARADDR_in_MD_CL1     ( data_master_CL1.ar_addr  ),
     .ARLEN_in_MD_CL1      ( data_master_CL1.ar_len   ),
     .ARSIZE_in_MD_CL1     ( data_master_CL1.ar_size  ),
     .ARBURST_in_MD_CL1    ( data_master_CL1.ar_burst ),
     .ARLOCK_in_MD_CL1     ( data_master_CL1.ar_lock  ),
     .ARCACHE_in_MD_CL1    ( data_master_CL1.ar_cache ),
     .ARPROT_in_MD_CL1     ( data_master_CL1.ar_prot  ),
     .ARVALID_in_MD_CL1    ( data_master_CL1.ar_valid ),
     .ARREADY_out_MD_CL1   ( data_master_CL1.ar_ready ),
     .RID_out_MD_CL1       ( data_master_CL1.r_id     ),
     .RDATA_out_MD_CL1     ( data_master_CL1.r_data   ),
     .RRESP_out_MD_CL1     ( data_master_CL1.r_resp   ),
     .RLAST_out_MD_CL1     ( data_master_CL1.r_last   ),
     .RVALID_out_MD_CL1    ( data_master_CL1.r_valid  ),
     .RREADY_in_MD_CL1     ( data_master_CL1.r_ready  ),
     .BID_out_MD_CL1       ( data_master_CL1.b_id     ),
     .BRESP_out_MD_CL1     ( data_master_CL1.b_resp   ),
     .BVALID_out_MD_CL1    ( data_master_CL1.b_valid  ),
     .BREADY_in_MD_CL1     ( data_master_CL1.b_ready  ),
     .init_div_MD_CL1      ( 1                        ),

     .AWID_in_MI_CL1       ( instr_master_CL1.aw_id    ),
     .AWADDR_in_MI_CL1     ( instr_master_CL1.aw_addr  ),
     .AWLEN_in_MI_CL1      ( instr_master_CL1.aw_len   ),
     .AWSIZE_in_MI_CL1     ( instr_master_CL1.aw_size  ),
     .AWBURST_in_MI_CL1    ( instr_master_CL1.aw_burst ),
     .AWLOCK_in_MI_CL1     ( instr_master_CL1.aw_lock  ),
     .AWCACHE_in_MI_CL1    ( instr_master_CL1.aw_cache ),
     .AWPROT_in_MI_CL1     ( instr_master_CL1.aw_prot  ),
     .AWVALID_in_MI_CL1    ( instr_master_CL1.aw_valid ),
     .AWREADY_out_MI_CL1   ( instr_master_CL1.aw_ready ),
     .WID_in_MI_CL1        ( '0                        ),
     .WDATA_in_MI_CL1      ( instr_master_CL1.w_data   ),
     .WSTRB_in_MI_CL1      ( instr_master_CL1.w_strb   ),
     .WLAST_in_MI_CL1      ( instr_master_CL1.w_last   ),
     .WVALID_in_MI_CL1     ( instr_master_CL1.w_valid  ),
     .WREADY_out_MI_CL1    ( instr_master_CL1.w_ready  ),
     .ARID_in_MI_CL1       ( instr_master_CL1.ar_id    ),
     .ARADDR_in_MI_CL1     ( instr_master_CL1.ar_addr  ),
     .ARLEN_in_MI_CL1      ( instr_master_CL1.ar_len   ),
     .ARSIZE_in_MI_CL1     ( instr_master_CL1.ar_size  ),
     .ARBURST_in_MI_CL1    ( instr_master_CL1.ar_burst ),
     .ARLOCK_in_MI_CL1     ( instr_master_CL1.ar_lock  ),
     .ARCACHE_in_MI_CL1    ( instr_master_CL1.ar_cache ),
     .ARPROT_in_MI_CL1     ( instr_master_CL1.ar_prot  ),
     .ARVALID_in_MI_CL1    ( instr_master_CL1.ar_valid ),
     .ARREADY_out_MI_CL1   ( instr_master_CL1.ar_ready ),
     .RID_out_MI_CL1       ( instr_master_CL1.r_id     ),
     .RDATA_out_MI_CL1     ( instr_master_CL1.r_data   ),
     .RRESP_out_MI_CL1     ( instr_master_CL1.r_resp   ),
     .RLAST_out_MI_CL1     ( instr_master_CL1.r_last   ),
     .RVALID_out_MI_CL1    ( instr_master_CL1.r_valid  ),
     .RREADY_in_MI_CL1     ( instr_master_CL1.r_ready  ),
     .BID_out_MI_CL1       ( instr_master_CL1.b_id     ),
     .BRESP_out_MI_CL1     ( instr_master_CL1.b_resp   ),
     .BVALID_out_MI_CL1    ( instr_master_CL1.b_valid  ),
     .BREADY_in_MI_CL1     ( instr_master_CL1.b_ready  ),
     .init_div_MI_CL1      ( 1                         ),

     .AWID_out_SD_CL1      ( data_slave_CL1.aw_id      ),
     .AWADDR_out_SD_CL1    ( data_slave_CL1.aw_addr    ),
     .AWLEN_out_SD_CL1     ( data_slave_CL1.aw_len     ),
     .AWSIZE_out_SD_CL1    ( data_slave_CL1.aw_size    ),
     .AWBURST_out_SD_CL1   ( data_slave_CL1.aw_burst   ),
     .AWLOCK_out_SD_CL1    ( data_slave_CL1.aw_lock    ),
     .AWCACHE_out_SD_CL1   ( data_slave_CL1.aw_cache   ),
     .AWPROT_out_SD_CL1    ( data_slave_CL1.aw_prot    ),
     .AWVALID_out_SD_CL1   ( data_slave_CL1.aw_valid   ),
     .AWREADY_in_SD_CL1    ( data_slave_CL1.aw_ready   ),
     .WID_out_SD_CL1       (                           ),
     .WDATA_out_SD_CL1     ( data_slave_CL1.w_data     ),
     .WSTRB_out_SD_CL1     ( data_slave_CL1.w_strb     ),
     .WLAST_out_SD_CL1     ( data_slave_CL1.w_last     ),
     .WVALID_out_SD_CL1    ( data_slave_CL1.w_valid    ),
     .WREADY_in_SD_CL1     ( data_slave_CL1.w_ready    ),
     .ARID_out_SD_CL1      ( data_slave_CL1.ar_id      ),
     .ARADDR_out_SD_CL1    ( data_slave_CL1.ar_addr    ),
     .ARLEN_out_SD_CL1     ( data_slave_CL1.ar_len     ),
     .ARSIZE_out_SD_CL1    ( data_slave_CL1.ar_size    ),
     .ARBURST_out_SD_CL1   ( data_slave_CL1.ar_burst   ),
     .ARLOCK_out_SD_CL1    ( data_slave_CL1.ar_lock    ),
     .ARCACHE_out_SD_CL1   ( data_slave_CL1.ar_cache   ),
     .ARPROT_out_SD_CL1    ( data_slave_CL1.ar_prot    ),
     .ARVALID_out_SD_CL1   ( data_slave_CL1.ar_valid   ),
     .ARREADY_in_SD_CL1    ( data_slave_CL1.ar_ready   ),
     .RID_in_SD_CL1        ( data_slave_CL1.r_id       ),
     .RDATA_in_SD_CL1      ( data_slave_CL1.r_data     ),
     .RRESP_in_SD_CL1      ( data_slave_CL1.r_resp     ),
     .RLAST_in_SD_CL1      ( data_slave_CL1.r_last     ),
     .RVALID_in_SD_CL1     ( data_slave_CL1.r_valid    ),
     .RREADY_out_SD_CL1    ( data_slave_CL1.r_ready    ),
     .BID_in_SD_CL1        ( data_slave_CL1.b_id       ),
     .BRESP_in_SD_CL1      ( data_slave_CL1.b_resp     ),
     .BVALID_in_SD_CL1     ( data_slave_CL1.b_valid    ),
     .BREADY_out_SD_CL1    ( data_slave_CL1.b_ready    ),
     .target_div_SD_CL1    ( 1                         ),

     .AWID_in_MD_CL2       ( data_master_CL2.aw_id     ),
     .AWADDR_in_MD_CL2     ( data_master_CL2.aw_addr   ),
     .AWLEN_in_MD_CL2      ( data_master_CL2.aw_len    ),
     .AWSIZE_in_MD_CL2     ( data_master_CL2.aw_size   ),
     .AWBURST_in_MD_CL2    ( data_master_CL2.aw_burst  ),
     .AWLOCK_in_MD_CL2     ( data_master_CL2.aw_lock   ),
     .AWCACHE_in_MD_CL2    ( data_master_CL2.aw_cache  ),
     .AWPROT_in_MD_CL2     ( data_master_CL2.aw_prot   ),
     .AWVALID_in_MD_CL2    ( data_master_CL2.aw_valid  ),
     .AWREADY_out_MD_CL2   ( data_master_CL2.aw_ready  ),
     .WID_in_MD_CL2        ( '0                        ),
     .WDATA_in_MD_CL2      ( data_master_CL2.w_data    ),
     .WSTRB_in_MD_CL2      ( data_master_CL2.w_strb    ),
     .WLAST_in_MD_CL2      ( data_master_CL2.w_last    ),
     .WVALID_in_MD_CL2     ( data_master_CL2.w_valid   ),
     .WREADY_out_MD_CL2    ( data_master_CL2.w_ready   ),
     .ARID_in_MD_CL2       ( data_master_CL2.ar_id     ),
     .ARADDR_in_MD_CL2     ( data_master_CL2.ar_addr   ),
     .ARLEN_in_MD_CL2      ( data_master_CL2.ar_len    ),
     .ARSIZE_in_MD_CL2     ( data_master_CL2.ar_size   ),
     .ARBURST_in_MD_CL2    ( data_master_CL2.ar_burst  ),
     .ARLOCK_in_MD_CL2     ( data_master_CL2.ar_lock   ),
     .ARCACHE_in_MD_CL2    ( data_master_CL2.ar_cache  ),
     .ARPROT_in_MD_CL2     ( data_master_CL2.ar_prot   ),
     .ARVALID_in_MD_CL2    ( data_master_CL2.ar_valid  ),
     .ARREADY_out_MD_CL2   ( data_master_CL2.ar_ready  ),
     .RID_out_MD_CL2       ( data_master_CL2.r_id      ),
     .RDATA_out_MD_CL2     ( data_master_CL2.r_data    ),
     .RRESP_out_MD_CL2     ( data_master_CL2.r_resp    ),
     .RLAST_out_MD_CL2     ( data_master_CL2.r_last    ),
     .RVALID_out_MD_CL2    ( data_master_CL2.r_valid   ),
     .RREADY_in_MD_CL2     ( data_master_CL2.r_ready   ),
     .BID_out_MD_CL2       ( data_master_CL2.b_id      ),
     .BRESP_out_MD_CL2     ( data_master_CL2.b_resp    ),
     .BVALID_out_MD_CL2    ( data_master_CL2.b_valid   ),
     .BREADY_in_MD_CL2     ( data_master_CL2.b_ready   ),
     .init_div_MD_CL2      ( 1                         ),

     .AWID_in_MI_CL2       ( instr_master_CL2.aw_id    ),
     .AWADDR_in_MI_CL2     ( instr_master_CL2.aw_addr  ),
     .AWLEN_in_MI_CL2      ( instr_master_CL2.aw_len   ),
     .AWSIZE_in_MI_CL2     ( instr_master_CL2.aw_size  ),
     .AWBURST_in_MI_CL2    ( instr_master_CL2.aw_burst ),
     .AWLOCK_in_MI_CL2     ( instr_master_CL2.aw_lock  ),
     .AWCACHE_in_MI_CL2    ( instr_master_CL2.aw_cache ),
     .AWPROT_in_MI_CL2     ( instr_master_CL2.aw_prot  ),
     .AWVALID_in_MI_CL2    ( instr_master_CL2.aw_valid ),
     .AWREADY_out_MI_CL2   ( instr_master_CL2.aw_ready ),
     .WID_in_MI_CL2        ( '0                        ),
     .WDATA_in_MI_CL2      ( instr_master_CL2.w_data   ),
     .WSTRB_in_MI_CL2      ( instr_master_CL2.w_strb   ),
     .WLAST_in_MI_CL2      ( instr_master_CL2.w_last   ),
     .WVALID_in_MI_CL2     ( instr_master_CL2.w_valid  ),
     .WREADY_out_MI_CL2    ( instr_master_CL2.w_ready  ),
     .ARID_in_MI_CL2       ( instr_master_CL2.ar_id    ),
     .ARADDR_in_MI_CL2     ( instr_master_CL2.ar_addr  ),
     .ARLEN_in_MI_CL2      ( instr_master_CL2.ar_len   ),
     .ARSIZE_in_MI_CL2     ( instr_master_CL2.ar_size  ),
     .ARBURST_in_MI_CL2    ( instr_master_CL2.ar_burst ),
     .ARLOCK_in_MI_CL2     ( instr_master_CL2.ar_lock  ),
     .ARCACHE_in_MI_CL2    ( instr_master_CL2.ar_cache ),
     .ARPROT_in_MI_CL2     ( instr_master_CL2.ar_prot  ),
     .ARVALID_in_MI_CL2    ( instr_master_CL2.ar_valid ),
     .ARREADY_out_MI_CL2   ( instr_master_CL2.ar_ready ),
     .RID_out_MI_CL2       ( instr_master_CL2.r_id     ),
     .RDATA_out_MI_CL2     ( instr_master_CL2.r_data   ),
     .RRESP_out_MI_CL2     ( instr_master_CL2.r_resp   ),
     .RLAST_out_MI_CL2     ( instr_master_CL2.r_last   ),
     .RVALID_out_MI_CL2    ( instr_master_CL2.r_valid  ),
     .RREADY_in_MI_CL2     ( instr_master_CL2.r_ready  ),
     .BID_out_MI_CL2       ( instr_master_CL2.b_id     ),
     .BRESP_out_MI_CL2     ( instr_master_CL2.b_resp   ),
     .BVALID_out_MI_CL2    ( instr_master_CL2.b_valid  ),
     .BREADY_in_MI_CL2     ( instr_master_CL2.b_ready  ),
     .init_div_MI_CL2      ( 1                         ),

     .AWID_out_SD_CL2      ( data_slave_CL2.aw_id      ),
     .AWADDR_out_SD_CL2    ( data_slave_CL2.aw_addr    ),
     .AWLEN_out_SD_CL2     ( data_slave_CL2.aw_len     ),
     .AWSIZE_out_SD_CL2    ( data_slave_CL2.aw_size    ),
     .AWBURST_out_SD_CL2   ( data_slave_CL2.aw_burst   ),
     .AWLOCK_out_SD_CL2    ( data_slave_CL2.aw_lock    ),
     .AWCACHE_out_SD_CL2   ( data_slave_CL2.aw_cache   ),
     .AWPROT_out_SD_CL2    ( data_slave_CL2.aw_prot    ),
     .AWVALID_out_SD_CL2   ( data_slave_CL2.aw_valid   ),
     .AWREADY_in_SD_CL2    ( data_slave_CL2.aw_ready   ),
     .WID_out_SD_CL2       (                           ),
     .WDATA_out_SD_CL2     ( data_slave_CL2.w_data     ),
     .WSTRB_out_SD_CL2     ( data_slave_CL2.w_strb     ),
     .WLAST_out_SD_CL2     ( data_slave_CL2.w_last     ),
     .WVALID_out_SD_CL2    ( data_slave_CL2.w_valid    ),
     .WREADY_in_SD_CL2     ( data_slave_CL2.w_ready    ),
     .ARID_out_SD_CL2      ( data_slave_CL2.ar_id      ),
     .ARADDR_out_SD_CL2    ( data_slave_CL2.ar_addr    ),
     .ARLEN_out_SD_CL2     ( data_slave_CL2.ar_len     ),
     .ARSIZE_out_SD_CL2    ( data_slave_CL2.ar_size    ),
     .ARBURST_out_SD_CL2   ( data_slave_CL2.ar_burst   ),
     .ARLOCK_out_SD_CL2    ( data_slave_CL2.ar_lock    ),
     .ARCACHE_out_SD_CL2   ( data_slave_CL2.ar_cache   ),
     .ARPROT_out_SD_CL2    ( data_slave_CL2.ar_prot    ),
     .ARVALID_out_SD_CL2   ( data_slave_CL2.ar_valid   ),
     .ARREADY_in_SD_CL2    ( data_slave_CL2.ar_ready   ),
     .RID_in_SD_CL2        ( data_slave_CL2.r_id       ),
     .RDATA_in_SD_CL2      ( data_slave_CL2.r_data     ),
     .RRESP_in_SD_CL2      ( data_slave_CL2.r_resp     ),
     .RLAST_in_SD_CL2      ( data_slave_CL2.r_last     ),
     .RVALID_in_SD_CL2     ( data_slave_CL2.r_valid    ),
     .RREADY_out_SD_CL2    ( data_slave_CL2.r_ready    ),
     .BID_in_SD_CL2        ( data_slave_CL2.b_id       ),
     .BRESP_in_SD_CL2      ( data_slave_CL2.b_resp     ),
     .BVALID_in_SD_CL2     ( data_slave_CL2.b_valid    ),
     .BREADY_out_SD_CL2    ( data_slave_CL2.b_ready    ),
     .target_div_SD_CL2    ( 1                         ),

     .AWID_in_MD_CL3       ( data_master_CL3.aw_id    ),
     .AWADDR_in_MD_CL3     ( data_master_CL3.aw_addr  ),
     .AWLEN_in_MD_CL3      ( data_master_CL3.aw_len   ),
     .AWSIZE_in_MD_CL3     ( data_master_CL3.aw_size  ),
     .AWBURST_in_MD_CL3    ( data_master_CL3.aw_burst ),
     .AWLOCK_in_MD_CL3     ( data_master_CL3.aw_lock  ),
     .AWCACHE_in_MD_CL3    ( data_master_CL3.aw_cache ),
     .AWPROT_in_MD_CL3     ( data_master_CL3.aw_prot  ),
     .AWVALID_in_MD_CL3    ( data_master_CL3.aw_valid ),
     .AWREADY_out_MD_CL3   ( data_master_CL3.aw_ready ),
     .WID_in_MD_CL3        ( '0                       ),
     .WDATA_in_MD_CL3      ( data_master_CL3.w_data   ),
     .WSTRB_in_MD_CL3      ( data_master_CL3.w_strb   ),
     .WLAST_in_MD_CL3      ( data_master_CL3.w_last   ),
     .WVALID_in_MD_CL3     ( data_master_CL3.w_valid  ),
     .WREADY_out_MD_CL3    ( data_master_CL3.w_ready  ),
     .ARID_in_MD_CL3       ( data_master_CL3.ar_id    ),
     .ARADDR_in_MD_CL3     ( data_master_CL3.ar_addr  ),
     .ARLEN_in_MD_CL3      ( data_master_CL3.ar_len   ),
     .ARSIZE_in_MD_CL3     ( data_master_CL3.ar_size  ),
     .ARBURST_in_MD_CL3    ( data_master_CL3.ar_burst ),
     .ARLOCK_in_MD_CL3     ( data_master_CL3.ar_lock  ),
     .ARCACHE_in_MD_CL3    ( data_master_CL3.ar_cache ),
     .ARPROT_in_MD_CL3     ( data_master_CL3.ar_prot  ),
     .ARVALID_in_MD_CL3    ( data_master_CL3.ar_valid ),
     .ARREADY_out_MD_CL3   ( data_master_CL3.ar_ready ),
     .RID_out_MD_CL3       ( data_master_CL3.r_id     ),
     .RDATA_out_MD_CL3     ( data_master_CL3.r_data   ),
     .RRESP_out_MD_CL3     ( data_master_CL3.r_resp   ),
     .RLAST_out_MD_CL3     ( data_master_CL3.r_last   ),
     .RVALID_out_MD_CL3    ( data_master_CL3.r_valid  ),
     .RREADY_in_MD_CL3     ( data_master_CL3.r_ready  ),
     .BID_out_MD_CL3       ( data_master_CL3.b_id     ),
     .BRESP_out_MD_CL3     ( data_master_CL3.b_resp   ),
     .BVALID_out_MD_CL3    ( data_master_CL3.b_valid  ),
     .BREADY_in_MD_CL3     ( data_master_CL3.b_ready  ),
     .init_div_MD_CL3      ( 1                        ),

     .AWID_in_MI_CL3       ( instr_master_CL3.aw_id    ),
     .AWADDR_in_MI_CL3     ( instr_master_CL3.aw_addr  ),
     .AWLEN_in_MI_CL3      ( instr_master_CL3.aw_len   ),
     .AWSIZE_in_MI_CL3     ( instr_master_CL3.aw_size  ),
     .AWBURST_in_MI_CL3    ( instr_master_CL3.aw_burst ),
     .AWLOCK_in_MI_CL3     ( instr_master_CL3.aw_lock  ),
     .AWCACHE_in_MI_CL3    ( instr_master_CL3.aw_cache ),
     .AWPROT_in_MI_CL3     ( instr_master_CL3.aw_prot  ),
     .AWVALID_in_MI_CL3    ( instr_master_CL3.aw_valid ),
     .AWREADY_out_MI_CL3   ( instr_master_CL3.aw_ready ),
     .WID_in_MI_CL3        ( '0                        ),
     .WDATA_in_MI_CL3      ( instr_master_CL3.w_data   ),
     .WSTRB_in_MI_CL3      ( instr_master_CL3.w_strb   ),
     .WLAST_in_MI_CL3      ( instr_master_CL3.w_last   ),
     .WVALID_in_MI_CL3     ( instr_master_CL3.w_valid  ),
     .WREADY_out_MI_CL3    ( instr_master_CL3.w_ready  ),
     .ARID_in_MI_CL3       ( instr_master_CL3.ar_id    ),
     .ARADDR_in_MI_CL3     ( instr_master_CL3.ar_addr  ),
     .ARLEN_in_MI_CL3      ( instr_master_CL3.ar_len   ),
     .ARSIZE_in_MI_CL3     ( instr_master_CL3.ar_size  ),
     .ARBURST_in_MI_CL3    ( instr_master_CL3.ar_burst ),
     .ARLOCK_in_MI_CL3     ( instr_master_CL3.ar_lock  ),
     .ARCACHE_in_MI_CL3    ( instr_master_CL3.ar_cache ),
     .ARPROT_in_MI_CL3     ( instr_master_CL3.ar_prot  ),
     .ARVALID_in_MI_CL3    ( instr_master_CL3.ar_valid ),
     .ARREADY_out_MI_CL3   ( instr_master_CL3.ar_ready ),
     .RID_out_MI_CL3       ( instr_master_CL3.r_id     ),
     .RDATA_out_MI_CL3     ( instr_master_CL3.r_data   ),
     .RRESP_out_MI_CL3     ( instr_master_CL3.r_resp   ),
     .RLAST_out_MI_CL3     ( instr_master_CL3.r_last   ),
     .RVALID_out_MI_CL3    ( instr_master_CL3.r_valid  ),
     .RREADY_in_MI_CL3     ( instr_master_CL3.r_ready  ),
     .BID_out_MI_CL3       ( instr_master_CL3.b_id     ),
     .BRESP_out_MI_CL3     ( instr_master_CL3.b_resp   ),
     .BVALID_out_MI_CL3    ( instr_master_CL3.b_valid  ),
     .BREADY_in_MI_CL3     ( instr_master_CL3.b_ready  ),
     .init_div_MI_CL3      ( 1                         ),

     .AWID_out_SD_CL3      ( data_slave_CL3.aw_id    ),
     .AWADDR_out_SD_CL3    ( data_slave_CL3.aw_addr  ),
     .AWLEN_out_SD_CL3     ( data_slave_CL3.aw_len   ),
     .AWSIZE_out_SD_CL3    ( data_slave_CL3.aw_size  ),
     .AWBURST_out_SD_CL3   ( data_slave_CL3.aw_burst ),
     .AWLOCK_out_SD_CL3    ( data_slave_CL3.aw_lock  ),
     .AWCACHE_out_SD_CL3   ( data_slave_CL3.aw_cache ),
     .AWPROT_out_SD_CL3    ( data_slave_CL3.aw_prot  ),
     .AWVALID_out_SD_CL3   ( data_slave_CL3.aw_valid ),
     .AWREADY_in_SD_CL3    ( data_slave_CL3.aw_ready ),
     .WID_out_SD_CL3       (                         ),
     .WDATA_out_SD_CL3     ( data_slave_CL3.w_data   ),
     .WSTRB_out_SD_CL3     ( data_slave_CL3.w_strb   ),
     .WLAST_out_SD_CL3     ( data_slave_CL3.w_last   ),
     .WVALID_out_SD_CL3    ( data_slave_CL3.w_valid  ),
     .WREADY_in_SD_CL3     ( data_slave_CL3.w_ready  ),
     .ARID_out_SD_CL3      ( data_slave_CL3.ar_id    ),
     .ARADDR_out_SD_CL3    ( data_slave_CL3.ar_addr  ),
     .ARLEN_out_SD_CL3     ( data_slave_CL3.ar_len   ),
     .ARSIZE_out_SD_CL3    ( data_slave_CL3.ar_size  ),
     .ARBURST_out_SD_CL3   ( data_slave_CL3.ar_burst ),
     .ARLOCK_out_SD_CL3    ( data_slave_CL3.ar_lock  ),
     .ARCACHE_out_SD_CL3   ( data_slave_CL3.ar_cache ),
     .ARPROT_out_SD_CL3    ( data_slave_CL3.ar_prot  ),
     .ARVALID_out_SD_CL3   ( data_slave_CL3.ar_valid ),
     .ARREADY_in_SD_CL3    ( data_slave_CL3.ar_ready ),
     .RID_in_SD_CL3        ( data_slave_CL3.r_id     ),
     .RDATA_in_SD_CL3      ( data_slave_CL3.r_data   ),
     .RRESP_in_SD_CL3      ( data_slave_CL3.r_resp   ),
     .RLAST_in_SD_CL3      ( data_slave_CL3.r_last   ),
     .RVALID_in_SD_CL3     ( data_slave_CL3.r_valid  ),
     .RREADY_out_SD_CL3    ( data_slave_CL3.r_ready  ),
     .BID_in_SD_CL3        ( data_slave_CL3.b_id     ),
     .BRESP_in_SD_CL3      ( data_slave_CL3.b_resp   ),
     .BVALID_in_SD_CL3     ( data_slave_CL3.b_valid  ),
     .BREADY_out_SD_CL3    ( data_slave_CL3.b_ready  ),
     .target_div_SD_CL3    ( 1                       ),

     .AWID_out_L2_MEM      ( data_master_L2_MEM.aw_id    ),
     .AWADDR_out_L2_MEM    ( data_master_L2_MEM.aw_addr  ),
     .AWLEN_out_L2_MEM     ( data_master_L2_MEM.aw_len   ),
     .AWSIZE_out_L2_MEM    ( data_master_L2_MEM.aw_size  ),
     .AWBURST_out_L2_MEM   ( data_master_L2_MEM.aw_burst ),
     .AWLOCK_out_L2_MEM    ( data_master_L2_MEM.aw_lock  ),
     .AWCACHE_out_L2_MEM   ( data_master_L2_MEM.aw_cache ),
     .AWPROT_out_L2_MEM    ( data_master_L2_MEM.aw_prot  ),
     .AWVALID_out_L2_MEM   ( data_master_L2_MEM.aw_valid ),
     .AWREADY_in_L2_MEM    ( data_master_L2_MEM.aw_ready ),
     .WID_out_L2_MEM       (                             ),
     .WDATA_out_L2_MEM     ( data_master_L2_MEM.w_data   ),
     .WSTRB_out_L2_MEM     ( data_master_L2_MEM.w_strb   ),
     .WLAST_out_L2_MEM     ( data_master_L2_MEM.w_last   ),
     .WVALID_out_L2_MEM    ( data_master_L2_MEM.w_valid  ),
     .WREADY_in_L2_MEM     ( data_master_L2_MEM.w_ready  ),
     .ARID_out_L2_MEM      ( data_master_L2_MEM.ar_id    ),
     .ARADDR_out_L2_MEM    ( data_master_L2_MEM.ar_addr  ),
     .ARLEN_out_L2_MEM     ( data_master_L2_MEM.ar_len   ),
     .ARSIZE_out_L2_MEM    ( data_master_L2_MEM.ar_size  ),
     .ARBURST_out_L2_MEM   ( data_master_L2_MEM.ar_burst ),
     .ARLOCK_out_L2_MEM    ( data_master_L2_MEM.ar_lock  ),
     .ARCACHE_out_L2_MEM   ( data_master_L2_MEM.ar_cache ),
     .ARPROT_out_L2_MEM    ( data_master_L2_MEM.ar_prot  ),
     .ARVALID_out_L2_MEM   ( data_master_L2_MEM.ar_valid ),
     .ARREADY_in_L2_MEM    ( data_master_L2_MEM.ar_ready ),
     .RID_in_L2_MEM        ( data_master_L2_MEM.r_id     ),
     .RDATA_in_L2_MEM      ( data_master_L2_MEM.r_data   ),
     .RRESP_in_L2_MEM      ( data_master_L2_MEM.r_resp   ),
     .RLAST_in_L2_MEM      ( data_master_L2_MEM.r_last   ),
     .RVALID_in_L2_MEM     ( data_master_L2_MEM.r_valid  ),
     .RREADY_out_L2_MEM    ( data_master_L2_MEM.r_ready  ),
     .BID_in_L2_MEM        ( data_master_L2_MEM.b_id     ),
     .BRESP_in_L2_MEM      ( data_master_L2_MEM.b_resp   ),
     .BVALID_in_L2_MEM     ( data_master_L2_MEM.b_valid  ),
     .BREADY_out_L2_MEM    ( data_master_L2_MEM.b_ready  ),
     .target_div_L2_MEM    ( 1                           ),

     .AWID_in_EXT          ( data_slave_EXT.aw_id    ),
     .AWADDR_in_EXT        ( data_slave_EXT.aw_addr  ),
     .AWLEN_in_EXT         ( data_slave_EXT.aw_len   ),
     .AWSIZE_in_EXT        ( data_slave_EXT.aw_size  ),
     .AWBURST_in_EXT       ( data_slave_EXT.aw_burst ),
     .AWLOCK_in_EXT        ( data_slave_EXT.aw_lock  ),
     .AWCACHE_in_EXT       ( data_slave_EXT.aw_cache ),
     .AWPROT_in_EXT        ( data_slave_EXT.aw_prot  ),
     .AWVALID_in_EXT       ( data_slave_EXT.aw_valid ),
     .AWREADY_out_EXT      ( data_slave_EXT.aw_ready ),
     .WID_in_EXT           (  '0                     ),
     .WDATA_in_EXT         ( data_slave_EXT.w_data   ),
     .WSTRB_in_EXT         ( data_slave_EXT.w_strb   ),
     .WLAST_in_EXT         ( data_slave_EXT.w_last   ),
     .WVALID_in_EXT        ( data_slave_EXT.w_valid  ),
     .WREADY_out_EXT       ( data_slave_EXT.w_ready  ),
     .ARID_in_EXT          ( data_slave_EXT.ar_id    ),
     .ARADDR_in_EXT        ( data_slave_EXT.ar_addr  ),
     .ARLEN_in_EXT         ( data_slave_EXT.ar_len   ),
     .ARSIZE_in_EXT        ( data_slave_EXT.ar_size  ),
     .ARBURST_in_EXT       ( data_slave_EXT.ar_burst ),
     .ARLOCK_in_EXT        ( data_slave_EXT.ar_lock  ),
     .ARCACHE_in_EXT       ( data_slave_EXT.ar_cache ),
     .ARPROT_in_EXT        ( data_slave_EXT.ar_prot  ),
     .ARVALID_in_EXT       ( data_slave_EXT.ar_valid ),
     .ARREADY_out_EXT      ( data_slave_EXT.ar_ready ),
     .RID_out_EXT          ( data_slave_EXT.r_id     ),
     .RDATA_out_EXT        ( data_slave_EXT.r_data   ),
     .RRESP_out_EXT        ( data_slave_EXT.r_resp   ),
     .RLAST_out_EXT        ( data_slave_EXT.r_last   ),
     .RVALID_out_EXT       ( data_slave_EXT.r_valid  ),
     .RREADY_in_EXT        ( data_slave_EXT.r_ready  ),
     .BID_out_EXT          ( data_slave_EXT.b_id     ),
     .BRESP_out_EXT        ( data_slave_EXT.b_resp   ),
     .BVALID_out_EXT       ( data_slave_EXT.b_valid  ),
     .BREADY_in_EXT        ( data_slave_EXT.b_ready  ),
     .init_div_EXT         ( 1                       )
);



endmodule // noc_interconnect_wrap