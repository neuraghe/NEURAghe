task ddr_w1_readmem_8x8_ramloops;
  $readmemh("slm_files/ddr_w1_mem_cut0_0.slm", `DDR_W1_BRAM_RAMLOOP(0) );
  $readmemh("slm_files/ddr_w1_mem_cut1_0.slm", `DDR_W1_BRAM_RAMLOOP(1) );
  $readmemh("slm_files/ddr_w1_mem_cut2_0.slm", `DDR_W1_BRAM_RAMLOOP(2) );
  $readmemh("slm_files/ddr_w1_mem_cut3_0.slm", `DDR_W1_BRAM_RAMLOOP(3) );
  $readmemh("slm_files/ddr_w1_mem_cut4_0.slm", `DDR_W1_BRAM_RAMLOOP(4) );
  $readmemh("slm_files/ddr_w1_mem_cut5_0.slm", `DDR_W1_BRAM_RAMLOOP(5) );
  $readmemh("slm_files/ddr_w1_mem_cut6_0.slm", `DDR_W1_BRAM_RAMLOOP(6) );
  $readmemh("slm_files/ddr_w1_mem_cut7_0.slm", `DDR_W1_BRAM_RAMLOOP(7) );
  $readmemh("slm_files/ddr_w1_mem_cut0_1.slm", `DDR_W1_BRAM_RAMLOOP(8) );
  $readmemh("slm_files/ddr_w1_mem_cut1_1.slm", `DDR_W1_BRAM_RAMLOOP(9) );
  $readmemh("slm_files/ddr_w1_mem_cut2_1.slm", `DDR_W1_BRAM_RAMLOOP(10) );
  $readmemh("slm_files/ddr_w1_mem_cut3_1.slm", `DDR_W1_BRAM_RAMLOOP(11) );
  $readmemh("slm_files/ddr_w1_mem_cut4_1.slm", `DDR_W1_BRAM_RAMLOOP(12) );
  $readmemh("slm_files/ddr_w1_mem_cut5_1.slm", `DDR_W1_BRAM_RAMLOOP(13) );
  $readmemh("slm_files/ddr_w1_mem_cut6_1.slm", `DDR_W1_BRAM_RAMLOOP(14) );
  $readmemh("slm_files/ddr_w1_mem_cut7_1.slm", `DDR_W1_BRAM_RAMLOOP(15) );
  $readmemh("slm_files/ddr_w1_mem_cut0_2.slm", `DDR_W1_BRAM_RAMLOOP(16) );
  $readmemh("slm_files/ddr_w1_mem_cut1_2.slm", `DDR_W1_BRAM_RAMLOOP(17) );
  $readmemh("slm_files/ddr_w1_mem_cut2_2.slm", `DDR_W1_BRAM_RAMLOOP(18) );
  $readmemh("slm_files/ddr_w1_mem_cut3_2.slm", `DDR_W1_BRAM_RAMLOOP(19) );
  $readmemh("slm_files/ddr_w1_mem_cut4_2.slm", `DDR_W1_BRAM_RAMLOOP(20) );
  $readmemh("slm_files/ddr_w1_mem_cut5_2.slm", `DDR_W1_BRAM_RAMLOOP(21) );
  $readmemh("slm_files/ddr_w1_mem_cut6_2.slm", `DDR_W1_BRAM_RAMLOOP(22) );
  $readmemh("slm_files/ddr_w1_mem_cut7_2.slm", `DDR_W1_BRAM_RAMLOOP(23) );
  $readmemh("slm_files/ddr_w1_mem_cut0_3.slm", `DDR_W1_BRAM_RAMLOOP(24) );
  $readmemh("slm_files/ddr_w1_mem_cut1_3.slm", `DDR_W1_BRAM_RAMLOOP(25) );
  $readmemh("slm_files/ddr_w1_mem_cut2_3.slm", `DDR_W1_BRAM_RAMLOOP(26) );
  $readmemh("slm_files/ddr_w1_mem_cut3_3.slm", `DDR_W1_BRAM_RAMLOOP(27) );
  $readmemh("slm_files/ddr_w1_mem_cut4_3.slm", `DDR_W1_BRAM_RAMLOOP(28) );
  $readmemh("slm_files/ddr_w1_mem_cut5_3.slm", `DDR_W1_BRAM_RAMLOOP(29) );
  $readmemh("slm_files/ddr_w1_mem_cut6_3.slm", `DDR_W1_BRAM_RAMLOOP(30) );
  $readmemh("slm_files/ddr_w1_mem_cut7_3.slm", `DDR_W1_BRAM_RAMLOOP(31) );
  $readmemh("slm_files/ddr_w1_mem_cut0_4.slm", `DDR_W1_BRAM_RAMLOOP(32) );
  $readmemh("slm_files/ddr_w1_mem_cut1_4.slm", `DDR_W1_BRAM_RAMLOOP(33) );
  $readmemh("slm_files/ddr_w1_mem_cut2_4.slm", `DDR_W1_BRAM_RAMLOOP(34) );
  $readmemh("slm_files/ddr_w1_mem_cut3_4.slm", `DDR_W1_BRAM_RAMLOOP(35) );
  $readmemh("slm_files/ddr_w1_mem_cut4_4.slm", `DDR_W1_BRAM_RAMLOOP(36) );
  $readmemh("slm_files/ddr_w1_mem_cut5_4.slm", `DDR_W1_BRAM_RAMLOOP(37) );
  $readmemh("slm_files/ddr_w1_mem_cut6_4.slm", `DDR_W1_BRAM_RAMLOOP(38) );
  $readmemh("slm_files/ddr_w1_mem_cut7_4.slm", `DDR_W1_BRAM_RAMLOOP(39) );
  $readmemh("slm_files/ddr_w1_mem_cut0_5.slm", `DDR_W1_BRAM_RAMLOOP(40) );
  $readmemh("slm_files/ddr_w1_mem_cut1_5.slm", `DDR_W1_BRAM_RAMLOOP(41) );
  $readmemh("slm_files/ddr_w1_mem_cut2_5.slm", `DDR_W1_BRAM_RAMLOOP(42) );
  $readmemh("slm_files/ddr_w1_mem_cut3_5.slm", `DDR_W1_BRAM_RAMLOOP(43) );
  $readmemh("slm_files/ddr_w1_mem_cut4_5.slm", `DDR_W1_BRAM_RAMLOOP(44) );
  $readmemh("slm_files/ddr_w1_mem_cut5_5.slm", `DDR_W1_BRAM_RAMLOOP(45) );
  $readmemh("slm_files/ddr_w1_mem_cut6_5.slm", `DDR_W1_BRAM_RAMLOOP(46) );
  $readmemh("slm_files/ddr_w1_mem_cut7_5.slm", `DDR_W1_BRAM_RAMLOOP(47) );
  $readmemh("slm_files/ddr_w1_mem_cut0_6.slm", `DDR_W1_BRAM_RAMLOOP(48) );
  $readmemh("slm_files/ddr_w1_mem_cut1_6.slm", `DDR_W1_BRAM_RAMLOOP(49) );
  $readmemh("slm_files/ddr_w1_mem_cut2_6.slm", `DDR_W1_BRAM_RAMLOOP(50) );
  $readmemh("slm_files/ddr_w1_mem_cut3_6.slm", `DDR_W1_BRAM_RAMLOOP(51) );
  $readmemh("slm_files/ddr_w1_mem_cut4_6.slm", `DDR_W1_BRAM_RAMLOOP(52) );
  $readmemh("slm_files/ddr_w1_mem_cut5_6.slm", `DDR_W1_BRAM_RAMLOOP(53) );
  $readmemh("slm_files/ddr_w1_mem_cut6_6.slm", `DDR_W1_BRAM_RAMLOOP(54) );
  $readmemh("slm_files/ddr_w1_mem_cut7_6.slm", `DDR_W1_BRAM_RAMLOOP(55) );
  $readmemh("slm_files/ddr_w1_mem_cut0_7.slm", `DDR_W1_BRAM_RAMLOOP(56) );
  $readmemh("slm_files/ddr_w1_mem_cut1_7.slm", `DDR_W1_BRAM_RAMLOOP(57) );
  $readmemh("slm_files/ddr_w1_mem_cut2_7.slm", `DDR_W1_BRAM_RAMLOOP(58) );
  $readmemh("slm_files/ddr_w1_mem_cut3_7.slm", `DDR_W1_BRAM_RAMLOOP(59) );
  $readmemh("slm_files/ddr_w1_mem_cut4_7.slm", `DDR_W1_BRAM_RAMLOOP(60) );
  $readmemh("slm_files/ddr_w1_mem_cut5_7.slm", `DDR_W1_BRAM_RAMLOOP(61) );
  $readmemh("slm_files/ddr_w1_mem_cut6_7.slm", `DDR_W1_BRAM_RAMLOOP(62) );
  $readmemh("slm_files/ddr_w1_mem_cut7_7.slm", `DDR_W1_BRAM_RAMLOOP(63) );
endtask
