///////////////////////////////////////////////////////////////////////////////
// Copyright 2009 iNoCs                                                      //
//                                                                           //
// name         /home/chester/Desktop/prj/XPIPES_fresh/inocs/flow/rtl/verilog/noc_interconnect.v                                     //
// author       Federico Angiolini - angiolini@inocs.com                     //
// author       Antonio Pullini - pullini@inocs.com                          //
// info         Describes a NoC interconnect.  //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////
//                                                                           //
///////////////////////////////////////////////////////////////////////////////
//                    Automatically generated - don't edit                   //
//           File generated for topology: noc18_4sw_80bits_run0           //
///////////////////////////////////////////////////////////////////////////////

`include "noc_parameters.v"

module noc_interconnect(clk, rst, AWID_in_MD_CL0, AWADDR_in_MD_CL0, AWLEN_in_MD_CL0, AWSIZE_in_MD_CL0, AWBURST_in_MD_CL0, AWLOCK_in_MD_CL0, AWCACHE_in_MD_CL0, AWPROT_in_MD_CL0, AWVALID_in_MD_CL0, AWREADY_out_MD_CL0, WID_in_MD_CL0, WDATA_in_MD_CL0, WSTRB_in_MD_CL0, WLAST_in_MD_CL0, WVALID_in_MD_CL0, WREADY_out_MD_CL0, ARID_in_MD_CL0, ARADDR_in_MD_CL0, ARLEN_in_MD_CL0, ARSIZE_in_MD_CL0, ARBURST_in_MD_CL0, ARLOCK_in_MD_CL0, ARCACHE_in_MD_CL0, ARPROT_in_MD_CL0, ARVALID_in_MD_CL0, ARREADY_out_MD_CL0, RID_out_MD_CL0, RDATA_out_MD_CL0, RRESP_out_MD_CL0, RLAST_out_MD_CL0, RVALID_out_MD_CL0, RREADY_in_MD_CL0, BID_out_MD_CL0, BRESP_out_MD_CL0, BVALID_out_MD_CL0, BREADY_in_MD_CL0, init_div_MD_CL0, AWID_out_SD_CL0, AWADDR_out_SD_CL0, AWLEN_out_SD_CL0, AWSIZE_out_SD_CL0, AWBURST_out_SD_CL0, AWLOCK_out_SD_CL0, AWCACHE_out_SD_CL0, AWPROT_out_SD_CL0, AWVALID_out_SD_CL0, AWREADY_in_SD_CL0, WID_out_SD_CL0, WDATA_out_SD_CL0, WSTRB_out_SD_CL0, WLAST_out_SD_CL0, WVALID_out_SD_CL0, WREADY_in_SD_CL0, ARID_out_SD_CL0, ARADDR_out_SD_CL0, ARLEN_out_SD_CL0, ARSIZE_out_SD_CL0, ARBURST_out_SD_CL0, ARLOCK_out_SD_CL0, ARCACHE_out_SD_CL0, ARPROT_out_SD_CL0, ARVALID_out_SD_CL0, ARREADY_in_SD_CL0, RID_in_SD_CL0, RDATA_in_SD_CL0, RRESP_in_SD_CL0, RLAST_in_SD_CL0, RVALID_in_SD_CL0, RREADY_out_SD_CL0, BID_in_SD_CL0, BRESP_in_SD_CL0, BVALID_in_SD_CL0, BREADY_out_SD_CL0, target_div_SD_CL0, AWID_in_MI_CL0, AWADDR_in_MI_CL0, AWLEN_in_MI_CL0, AWSIZE_in_MI_CL0, AWBURST_in_MI_CL0, AWLOCK_in_MI_CL0, AWCACHE_in_MI_CL0, AWPROT_in_MI_CL0, AWVALID_in_MI_CL0, AWREADY_out_MI_CL0, WID_in_MI_CL0, WDATA_in_MI_CL0, WSTRB_in_MI_CL0, WLAST_in_MI_CL0, WVALID_in_MI_CL0, WREADY_out_MI_CL0, ARID_in_MI_CL0, ARADDR_in_MI_CL0, ARLEN_in_MI_CL0, ARSIZE_in_MI_CL0, ARBURST_in_MI_CL0, ARLOCK_in_MI_CL0, ARCACHE_in_MI_CL0, ARPROT_in_MI_CL0, ARVALID_in_MI_CL0, ARREADY_out_MI_CL0, RID_out_MI_CL0, RDATA_out_MI_CL0, RRESP_out_MI_CL0, RLAST_out_MI_CL0, RVALID_out_MI_CL0, RREADY_in_MI_CL0, BID_out_MI_CL0, BRESP_out_MI_CL0, BVALID_out_MI_CL0, BREADY_in_MI_CL0, init_div_MI_CL0, AWID_in_MD_CL1, AWADDR_in_MD_CL1, AWLEN_in_MD_CL1, AWSIZE_in_MD_CL1, AWBURST_in_MD_CL1, AWLOCK_in_MD_CL1, AWCACHE_in_MD_CL1, AWPROT_in_MD_CL1, AWVALID_in_MD_CL1, AWREADY_out_MD_CL1, WID_in_MD_CL1, WDATA_in_MD_CL1, WSTRB_in_MD_CL1, WLAST_in_MD_CL1, WVALID_in_MD_CL1, WREADY_out_MD_CL1, ARID_in_MD_CL1, ARADDR_in_MD_CL1, ARLEN_in_MD_CL1, ARSIZE_in_MD_CL1, ARBURST_in_MD_CL1, ARLOCK_in_MD_CL1, ARCACHE_in_MD_CL1, ARPROT_in_MD_CL1, ARVALID_in_MD_CL1, ARREADY_out_MD_CL1, RID_out_MD_CL1, RDATA_out_MD_CL1, RRESP_out_MD_CL1, RLAST_out_MD_CL1, RVALID_out_MD_CL1, RREADY_in_MD_CL1, BID_out_MD_CL1, BRESP_out_MD_CL1, BVALID_out_MD_CL1, BREADY_in_MD_CL1, init_div_MD_CL1, AWID_in_MI_CL1, AWADDR_in_MI_CL1, AWLEN_in_MI_CL1, AWSIZE_in_MI_CL1, AWBURST_in_MI_CL1, AWLOCK_in_MI_CL1, AWCACHE_in_MI_CL1, AWPROT_in_MI_CL1, AWVALID_in_MI_CL1, AWREADY_out_MI_CL1, WID_in_MI_CL1, WDATA_in_MI_CL1, WSTRB_in_MI_CL1, WLAST_in_MI_CL1, WVALID_in_MI_CL1, WREADY_out_MI_CL1, ARID_in_MI_CL1, ARADDR_in_MI_CL1, ARLEN_in_MI_CL1, ARSIZE_in_MI_CL1, ARBURST_in_MI_CL1, ARLOCK_in_MI_CL1, ARCACHE_in_MI_CL1, ARPROT_in_MI_CL1, ARVALID_in_MI_CL1, ARREADY_out_MI_CL1, RID_out_MI_CL1, RDATA_out_MI_CL1, RRESP_out_MI_CL1, RLAST_out_MI_CL1, RVALID_out_MI_CL1, RREADY_in_MI_CL1, BID_out_MI_CL1, BRESP_out_MI_CL1, BVALID_out_MI_CL1, BREADY_in_MI_CL1, init_div_MI_CL1, AWID_out_SD_CL1, AWADDR_out_SD_CL1, AWLEN_out_SD_CL1, AWSIZE_out_SD_CL1, AWBURST_out_SD_CL1, AWLOCK_out_SD_CL1, AWCACHE_out_SD_CL1, AWPROT_out_SD_CL1, AWVALID_out_SD_CL1, AWREADY_in_SD_CL1, WID_out_SD_CL1, WDATA_out_SD_CL1, WSTRB_out_SD_CL1, WLAST_out_SD_CL1, WVALID_out_SD_CL1, WREADY_in_SD_CL1, ARID_out_SD_CL1, ARADDR_out_SD_CL1, ARLEN_out_SD_CL1, ARSIZE_out_SD_CL1, ARBURST_out_SD_CL1, ARLOCK_out_SD_CL1, ARCACHE_out_SD_CL1, ARPROT_out_SD_CL1, ARVALID_out_SD_CL1, ARREADY_in_SD_CL1, RID_in_SD_CL1, RDATA_in_SD_CL1, RRESP_in_SD_CL1, RLAST_in_SD_CL1, RVALID_in_SD_CL1, RREADY_out_SD_CL1, BID_in_SD_CL1, BRESP_in_SD_CL1, BVALID_in_SD_CL1, BREADY_out_SD_CL1, target_div_SD_CL1, AWID_in_MD_CL2, AWADDR_in_MD_CL2, AWLEN_in_MD_CL2, AWSIZE_in_MD_CL2, AWBURST_in_MD_CL2, AWLOCK_in_MD_CL2, AWCACHE_in_MD_CL2, AWPROT_in_MD_CL2, AWVALID_in_MD_CL2, AWREADY_out_MD_CL2, WID_in_MD_CL2, WDATA_in_MD_CL2, WSTRB_in_MD_CL2, WLAST_in_MD_CL2, WVALID_in_MD_CL2, WREADY_out_MD_CL2, ARID_in_MD_CL2, ARADDR_in_MD_CL2, ARLEN_in_MD_CL2, ARSIZE_in_MD_CL2, ARBURST_in_MD_CL2, ARLOCK_in_MD_CL2, ARCACHE_in_MD_CL2, ARPROT_in_MD_CL2, ARVALID_in_MD_CL2, ARREADY_out_MD_CL2, RID_out_MD_CL2, RDATA_out_MD_CL2, RRESP_out_MD_CL2, RLAST_out_MD_CL2, RVALID_out_MD_CL2, RREADY_in_MD_CL2, BID_out_MD_CL2, BRESP_out_MD_CL2, BVALID_out_MD_CL2, BREADY_in_MD_CL2, init_div_MD_CL2, AWID_in_MI_CL2, AWADDR_in_MI_CL2, AWLEN_in_MI_CL2, AWSIZE_in_MI_CL2, AWBURST_in_MI_CL2, AWLOCK_in_MI_CL2, AWCACHE_in_MI_CL2, AWPROT_in_MI_CL2, AWVALID_in_MI_CL2, AWREADY_out_MI_CL2, WID_in_MI_CL2, WDATA_in_MI_CL2, WSTRB_in_MI_CL2, WLAST_in_MI_CL2, WVALID_in_MI_CL2, WREADY_out_MI_CL2, ARID_in_MI_CL2, ARADDR_in_MI_CL2, ARLEN_in_MI_CL2, ARSIZE_in_MI_CL2, ARBURST_in_MI_CL2, ARLOCK_in_MI_CL2, ARCACHE_in_MI_CL2, ARPROT_in_MI_CL2, ARVALID_in_MI_CL2, ARREADY_out_MI_CL2, RID_out_MI_CL2, RDATA_out_MI_CL2, RRESP_out_MI_CL2, RLAST_out_MI_CL2, RVALID_out_MI_CL2, RREADY_in_MI_CL2, BID_out_MI_CL2, BRESP_out_MI_CL2, BVALID_out_MI_CL2, BREADY_in_MI_CL2, init_div_MI_CL2, AWID_out_SD_CL2, AWADDR_out_SD_CL2, AWLEN_out_SD_CL2, AWSIZE_out_SD_CL2, AWBURST_out_SD_CL2, AWLOCK_out_SD_CL2, AWCACHE_out_SD_CL2, AWPROT_out_SD_CL2, AWVALID_out_SD_CL2, AWREADY_in_SD_CL2, WID_out_SD_CL2, WDATA_out_SD_CL2, WSTRB_out_SD_CL2, WLAST_out_SD_CL2, WVALID_out_SD_CL2, WREADY_in_SD_CL2, ARID_out_SD_CL2, ARADDR_out_SD_CL2, ARLEN_out_SD_CL2, ARSIZE_out_SD_CL2, ARBURST_out_SD_CL2, ARLOCK_out_SD_CL2, ARCACHE_out_SD_CL2, ARPROT_out_SD_CL2, ARVALID_out_SD_CL2, ARREADY_in_SD_CL2, RID_in_SD_CL2, RDATA_in_SD_CL2, RRESP_in_SD_CL2, RLAST_in_SD_CL2, RVALID_in_SD_CL2, RREADY_out_SD_CL2, BID_in_SD_CL2, BRESP_in_SD_CL2, BVALID_in_SD_CL2, BREADY_out_SD_CL2, target_div_SD_CL2, AWID_in_MD_CL3, AWADDR_in_MD_CL3, AWLEN_in_MD_CL3, AWSIZE_in_MD_CL3, AWBURST_in_MD_CL3, AWLOCK_in_MD_CL3, AWCACHE_in_MD_CL3, AWPROT_in_MD_CL3, AWVALID_in_MD_CL3, AWREADY_out_MD_CL3, WID_in_MD_CL3, WDATA_in_MD_CL3, WSTRB_in_MD_CL3, WLAST_in_MD_CL3, WVALID_in_MD_CL3, WREADY_out_MD_CL3, ARID_in_MD_CL3, ARADDR_in_MD_CL3, ARLEN_in_MD_CL3, ARSIZE_in_MD_CL3, ARBURST_in_MD_CL3, ARLOCK_in_MD_CL3, ARCACHE_in_MD_CL3, ARPROT_in_MD_CL3, ARVALID_in_MD_CL3, ARREADY_out_MD_CL3, RID_out_MD_CL3, RDATA_out_MD_CL3, RRESP_out_MD_CL3, RLAST_out_MD_CL3, RVALID_out_MD_CL3, RREADY_in_MD_CL3, BID_out_MD_CL3, BRESP_out_MD_CL3, BVALID_out_MD_CL3, BREADY_in_MD_CL3, init_div_MD_CL3, AWID_in_MI_CL3, AWADDR_in_MI_CL3, AWLEN_in_MI_CL3, AWSIZE_in_MI_CL3, AWBURST_in_MI_CL3, AWLOCK_in_MI_CL3, AWCACHE_in_MI_CL3, AWPROT_in_MI_CL3, AWVALID_in_MI_CL3, AWREADY_out_MI_CL3, WID_in_MI_CL3, WDATA_in_MI_CL3, WSTRB_in_MI_CL3, WLAST_in_MI_CL3, WVALID_in_MI_CL3, WREADY_out_MI_CL3, ARID_in_MI_CL3, ARADDR_in_MI_CL3, ARLEN_in_MI_CL3, ARSIZE_in_MI_CL3, ARBURST_in_MI_CL3, ARLOCK_in_MI_CL3, ARCACHE_in_MI_CL3, ARPROT_in_MI_CL3, ARVALID_in_MI_CL3, ARREADY_out_MI_CL3, RID_out_MI_CL3, RDATA_out_MI_CL3, RRESP_out_MI_CL3, RLAST_out_MI_CL3, RVALID_out_MI_CL3, RREADY_in_MI_CL3, BID_out_MI_CL3, BRESP_out_MI_CL3, BVALID_out_MI_CL3, BREADY_in_MI_CL3, init_div_MI_CL3, AWID_out_SD_CL3, AWADDR_out_SD_CL3, AWLEN_out_SD_CL3, AWSIZE_out_SD_CL3, AWBURST_out_SD_CL3, AWLOCK_out_SD_CL3, AWCACHE_out_SD_CL3, AWPROT_out_SD_CL3, AWVALID_out_SD_CL3, AWREADY_in_SD_CL3, WID_out_SD_CL3, WDATA_out_SD_CL3, WSTRB_out_SD_CL3, WLAST_out_SD_CL3, WVALID_out_SD_CL3, WREADY_in_SD_CL3, ARID_out_SD_CL3, ARADDR_out_SD_CL3, ARLEN_out_SD_CL3, ARSIZE_out_SD_CL3, ARBURST_out_SD_CL3, ARLOCK_out_SD_CL3, ARCACHE_out_SD_CL3, ARPROT_out_SD_CL3, ARVALID_out_SD_CL3, ARREADY_in_SD_CL3, RID_in_SD_CL3, RDATA_in_SD_CL3, RRESP_in_SD_CL3, RLAST_in_SD_CL3, RVALID_in_SD_CL3, RREADY_out_SD_CL3, BID_in_SD_CL3, BRESP_in_SD_CL3, BVALID_in_SD_CL3, BREADY_out_SD_CL3, target_div_SD_CL3, AWID_out_L2_MEM, AWADDR_out_L2_MEM, AWLEN_out_L2_MEM, AWSIZE_out_L2_MEM, AWBURST_out_L2_MEM, AWLOCK_out_L2_MEM, AWCACHE_out_L2_MEM, AWPROT_out_L2_MEM, AWVALID_out_L2_MEM, AWREADY_in_L2_MEM, WID_out_L2_MEM, WDATA_out_L2_MEM, WSTRB_out_L2_MEM, WLAST_out_L2_MEM, WVALID_out_L2_MEM, WREADY_in_L2_MEM, ARID_out_L2_MEM, ARADDR_out_L2_MEM, ARLEN_out_L2_MEM, ARSIZE_out_L2_MEM, ARBURST_out_L2_MEM, ARLOCK_out_L2_MEM, ARCACHE_out_L2_MEM, ARPROT_out_L2_MEM, ARVALID_out_L2_MEM, ARREADY_in_L2_MEM, RID_in_L2_MEM, RDATA_in_L2_MEM, RRESP_in_L2_MEM, RLAST_in_L2_MEM, RVALID_in_L2_MEM, RREADY_out_L2_MEM, BID_in_L2_MEM, BRESP_in_L2_MEM, BVALID_in_L2_MEM, BREADY_out_L2_MEM, target_div_L2_MEM, AWID_in_EXT, AWADDR_in_EXT, AWLEN_in_EXT, AWSIZE_in_EXT, AWBURST_in_EXT, AWLOCK_in_EXT, AWCACHE_in_EXT, AWPROT_in_EXT, AWVALID_in_EXT, AWREADY_out_EXT, WID_in_EXT, WDATA_in_EXT, WSTRB_in_EXT, WLAST_in_EXT, WVALID_in_EXT, WREADY_out_EXT, ARID_in_EXT, ARADDR_in_EXT, ARLEN_in_EXT, ARSIZE_in_EXT, ARBURST_in_EXT, ARLOCK_in_EXT, ARCACHE_in_EXT, ARPROT_in_EXT, ARVALID_in_EXT, ARREADY_out_EXT, RID_out_EXT, RDATA_out_EXT, RRESP_out_EXT, RLAST_out_EXT, RVALID_out_EXT, RREADY_in_EXT, BID_out_EXT, BRESP_out_EXT, BVALID_out_EXT, BREADY_in_EXT, init_div_EXT);

    input rst;
    input clk;
    input [3 : 0]                   AWID_in_MD_CL0;
    input [31 : 0]                  AWADDR_in_MD_CL0;
    input [7 : 0]                   AWLEN_in_MD_CL0;
    input [2 : 0]                   AWSIZE_in_MD_CL0;
    input [1 : 0]                   AWBURST_in_MD_CL0;
    input [1 : 0]                   AWLOCK_in_MD_CL0;
    input [3 : 0]                   AWCACHE_in_MD_CL0;
    input [2 : 0]                   AWPROT_in_MD_CL0;
    input                           AWVALID_in_MD_CL0;
    output                          AWREADY_out_MD_CL0;
    input [3 : 0]                   WID_in_MD_CL0;
    input [63 : 0]                  WDATA_in_MD_CL0;
    input [7 : 0]                   WSTRB_in_MD_CL0;
    input                           WLAST_in_MD_CL0;
    input                           WVALID_in_MD_CL0;
    output                          WREADY_out_MD_CL0;
    output [3 : 0]                  BID_out_MD_CL0;
    output [1 : 0]                  BRESP_out_MD_CL0;
    output                          BVALID_out_MD_CL0;
    input                           BREADY_in_MD_CL0;
    input [3 : 0]                   ARID_in_MD_CL0;
    input [31 : 0]                  ARADDR_in_MD_CL0;
    input [7 : 0]                   ARLEN_in_MD_CL0;
    input [2 : 0]                   ARSIZE_in_MD_CL0;
    input [1 : 0]                   ARBURST_in_MD_CL0;
    input [1 : 0]                   ARLOCK_in_MD_CL0;
    input [3 : 0]                   ARCACHE_in_MD_CL0;
    input [2 : 0]                   ARPROT_in_MD_CL0;
    input                           ARVALID_in_MD_CL0;
    output                          ARREADY_out_MD_CL0;
    output [3 : 0]                  RID_out_MD_CL0;
    output [63 : 0]                 RDATA_out_MD_CL0;
    output [1 : 0]                  RRESP_out_MD_CL0;
    output                          RLAST_out_MD_CL0;
    output                          RVALID_out_MD_CL0;
    input                           RREADY_in_MD_CL0;
    input [`COUNTERWD - 1 : 0]      init_div_MD_CL0;
    output [3 : 0]                  AWID_out_SD_CL0;
    output [31 : 0]                 AWADDR_out_SD_CL0;
    output [7 : 0]                  AWLEN_out_SD_CL0;
    output [2 : 0]                  AWSIZE_out_SD_CL0;
    output [1 : 0]                  AWBURST_out_SD_CL0;
    output [1 : 0]                  AWLOCK_out_SD_CL0;
    output [3 : 0]                  AWCACHE_out_SD_CL0;
    output [2 : 0]                  AWPROT_out_SD_CL0;
    output                          AWVALID_out_SD_CL0;
    input                           AWREADY_in_SD_CL0;
    output [3 : 0]                  WID_out_SD_CL0;
    output [63 : 0]                 WDATA_out_SD_CL0;
    output [7 : 0]                  WSTRB_out_SD_CL0;
    output                          WLAST_out_SD_CL0;
    output                          WVALID_out_SD_CL0;
    input                           WREADY_in_SD_CL0;
    input [3 : 0]                   BID_in_SD_CL0;
    input [1 : 0]                   BRESP_in_SD_CL0;
    input                           BVALID_in_SD_CL0;
    output                          BREADY_out_SD_CL0;
    output [3 : 0]                  ARID_out_SD_CL0;
    output [31 : 0]                 ARADDR_out_SD_CL0;
    output [7 : 0]                  ARLEN_out_SD_CL0;
    output [2 : 0]                  ARSIZE_out_SD_CL0;
    output [1 : 0]                  ARBURST_out_SD_CL0;
    output [1 : 0]                  ARLOCK_out_SD_CL0;
    output [3 : 0]                  ARCACHE_out_SD_CL0;
    output [2 : 0]                  ARPROT_out_SD_CL0;
    output                          ARVALID_out_SD_CL0;
    input                           ARREADY_in_SD_CL0;
    input [3 : 0]                   RID_in_SD_CL0;
    input [63 : 0]                  RDATA_in_SD_CL0;
    input [1 : 0]                   RRESP_in_SD_CL0;
    input                           RLAST_in_SD_CL0;
    input                           RVALID_in_SD_CL0;
    output                          RREADY_out_SD_CL0;
    input [`COUNTERWD - 1 : 0]      target_div_SD_CL0;
    input [3 : 0]                   AWID_in_MI_CL0;
    input [31 : 0]                  AWADDR_in_MI_CL0;
    input [7 : 0]                   AWLEN_in_MI_CL0;
    input [2 : 0]                   AWSIZE_in_MI_CL0;
    input [1 : 0]                   AWBURST_in_MI_CL0;
    input [1 : 0]                   AWLOCK_in_MI_CL0;
    input [3 : 0]                   AWCACHE_in_MI_CL0;
    input [2 : 0]                   AWPROT_in_MI_CL0;
    input                           AWVALID_in_MI_CL0;
    output                          AWREADY_out_MI_CL0;
    input [3 : 0]                   WID_in_MI_CL0;
    input [63 : 0]                  WDATA_in_MI_CL0;
    input [7 : 0]                   WSTRB_in_MI_CL0;
    input                           WLAST_in_MI_CL0;
    input                           WVALID_in_MI_CL0;
    output                          WREADY_out_MI_CL0;
    output [3 : 0]                  BID_out_MI_CL0;
    output [1 : 0]                  BRESP_out_MI_CL0;
    output                          BVALID_out_MI_CL0;
    input                           BREADY_in_MI_CL0;
    input [3 : 0]                   ARID_in_MI_CL0;
    input [31 : 0]                  ARADDR_in_MI_CL0;
    input [7 : 0]                   ARLEN_in_MI_CL0;
    input [2 : 0]                   ARSIZE_in_MI_CL0;
    input [1 : 0]                   ARBURST_in_MI_CL0;
    input [1 : 0]                   ARLOCK_in_MI_CL0;
    input [3 : 0]                   ARCACHE_in_MI_CL0;
    input [2 : 0]                   ARPROT_in_MI_CL0;
    input                           ARVALID_in_MI_CL0;
    output                          ARREADY_out_MI_CL0;
    output [3 : 0]                  RID_out_MI_CL0;
    output [63 : 0]                 RDATA_out_MI_CL0;
    output [1 : 0]                  RRESP_out_MI_CL0;
    output                          RLAST_out_MI_CL0;
    output                          RVALID_out_MI_CL0;
    input                           RREADY_in_MI_CL0;
    input [`COUNTERWD - 1 : 0]      init_div_MI_CL0;
    input [3 : 0]                   AWID_in_MD_CL1;
    input [31 : 0]                  AWADDR_in_MD_CL1;
    input [7 : 0]                   AWLEN_in_MD_CL1;
    input [2 : 0]                   AWSIZE_in_MD_CL1;
    input [1 : 0]                   AWBURST_in_MD_CL1;
    input [1 : 0]                   AWLOCK_in_MD_CL1;
    input [3 : 0]                   AWCACHE_in_MD_CL1;
    input [2 : 0]                   AWPROT_in_MD_CL1;
    input                           AWVALID_in_MD_CL1;
    output                          AWREADY_out_MD_CL1;
    input [3 : 0]                   WID_in_MD_CL1;
    input [63 : 0]                  WDATA_in_MD_CL1;
    input [7 : 0]                   WSTRB_in_MD_CL1;
    input                           WLAST_in_MD_CL1;
    input                           WVALID_in_MD_CL1;
    output                          WREADY_out_MD_CL1;
    output [3 : 0]                  BID_out_MD_CL1;
    output [1 : 0]                  BRESP_out_MD_CL1;
    output                          BVALID_out_MD_CL1;
    input                           BREADY_in_MD_CL1;
    input [3 : 0]                   ARID_in_MD_CL1;
    input [31 : 0]                  ARADDR_in_MD_CL1;
    input [7 : 0]                   ARLEN_in_MD_CL1;
    input [2 : 0]                   ARSIZE_in_MD_CL1;
    input [1 : 0]                   ARBURST_in_MD_CL1;
    input [1 : 0]                   ARLOCK_in_MD_CL1;
    input [3 : 0]                   ARCACHE_in_MD_CL1;
    input [2 : 0]                   ARPROT_in_MD_CL1;
    input                           ARVALID_in_MD_CL1;
    output                          ARREADY_out_MD_CL1;
    output [3 : 0]                  RID_out_MD_CL1;
    output [63 : 0]                 RDATA_out_MD_CL1;
    output [1 : 0]                  RRESP_out_MD_CL1;
    output                          RLAST_out_MD_CL1;
    output                          RVALID_out_MD_CL1;
    input                           RREADY_in_MD_CL1;
    input [`COUNTERWD - 1 : 0]      init_div_MD_CL1;
    input [3 : 0]                   AWID_in_MI_CL1;
    input [31 : 0]                  AWADDR_in_MI_CL1;
    input [7 : 0]                   AWLEN_in_MI_CL1;
    input [2 : 0]                   AWSIZE_in_MI_CL1;
    input [1 : 0]                   AWBURST_in_MI_CL1;
    input [1 : 0]                   AWLOCK_in_MI_CL1;
    input [3 : 0]                   AWCACHE_in_MI_CL1;
    input [2 : 0]                   AWPROT_in_MI_CL1;
    input                           AWVALID_in_MI_CL1;
    output                          AWREADY_out_MI_CL1;
    input [3 : 0]                   WID_in_MI_CL1;
    input [63 : 0]                  WDATA_in_MI_CL1;
    input [7 : 0]                   WSTRB_in_MI_CL1;
    input                           WLAST_in_MI_CL1;
    input                           WVALID_in_MI_CL1;
    output                          WREADY_out_MI_CL1;
    output [3 : 0]                  BID_out_MI_CL1;
    output [1 : 0]                  BRESP_out_MI_CL1;
    output                          BVALID_out_MI_CL1;
    input                           BREADY_in_MI_CL1;
    input [3 : 0]                   ARID_in_MI_CL1;
    input [31 : 0]                  ARADDR_in_MI_CL1;
    input [7 : 0]                   ARLEN_in_MI_CL1;
    input [2 : 0]                   ARSIZE_in_MI_CL1;
    input [1 : 0]                   ARBURST_in_MI_CL1;
    input [1 : 0]                   ARLOCK_in_MI_CL1;
    input [3 : 0]                   ARCACHE_in_MI_CL1;
    input [2 : 0]                   ARPROT_in_MI_CL1;
    input                           ARVALID_in_MI_CL1;
    output                          ARREADY_out_MI_CL1;
    output [3 : 0]                  RID_out_MI_CL1;
    output [63 : 0]                 RDATA_out_MI_CL1;
    output [1 : 0]                  RRESP_out_MI_CL1;
    output                          RLAST_out_MI_CL1;
    output                          RVALID_out_MI_CL1;
    input                           RREADY_in_MI_CL1;
    input [`COUNTERWD - 1 : 0]      init_div_MI_CL1;
    output [3 : 0]                  AWID_out_SD_CL1;
    output [31 : 0]                 AWADDR_out_SD_CL1;
    output [7 : 0]                  AWLEN_out_SD_CL1;
    output [2 : 0]                  AWSIZE_out_SD_CL1;
    output [1 : 0]                  AWBURST_out_SD_CL1;
    output [1 : 0]                  AWLOCK_out_SD_CL1;
    output [3 : 0]                  AWCACHE_out_SD_CL1;
    output [2 : 0]                  AWPROT_out_SD_CL1;
    output                          AWVALID_out_SD_CL1;
    input                           AWREADY_in_SD_CL1;
    output [3 : 0]                  WID_out_SD_CL1;
    output [63 : 0]                 WDATA_out_SD_CL1;
    output [7 : 0]                  WSTRB_out_SD_CL1;
    output                          WLAST_out_SD_CL1;
    output                          WVALID_out_SD_CL1;
    input                           WREADY_in_SD_CL1;
    input [3 : 0]                   BID_in_SD_CL1;
    input [1 : 0]                   BRESP_in_SD_CL1;
    input                           BVALID_in_SD_CL1;
    output                          BREADY_out_SD_CL1;
    output [3 : 0]                  ARID_out_SD_CL1;
    output [31 : 0]                 ARADDR_out_SD_CL1;
    output [7 : 0]                  ARLEN_out_SD_CL1;
    output [2 : 0]                  ARSIZE_out_SD_CL1;
    output [1 : 0]                  ARBURST_out_SD_CL1;
    output [1 : 0]                  ARLOCK_out_SD_CL1;
    output [3 : 0]                  ARCACHE_out_SD_CL1;
    output [2 : 0]                  ARPROT_out_SD_CL1;
    output                          ARVALID_out_SD_CL1;
    input                           ARREADY_in_SD_CL1;
    input [3 : 0]                   RID_in_SD_CL1;
    input [63 : 0]                  RDATA_in_SD_CL1;
    input [1 : 0]                   RRESP_in_SD_CL1;
    input                           RLAST_in_SD_CL1;
    input                           RVALID_in_SD_CL1;
    output                          RREADY_out_SD_CL1;
    input [`COUNTERWD - 1 : 0]      target_div_SD_CL1;
    input [3 : 0]                   AWID_in_MD_CL2;
    input [31 : 0]                  AWADDR_in_MD_CL2;
    input [7 : 0]                   AWLEN_in_MD_CL2;
    input [2 : 0]                   AWSIZE_in_MD_CL2;
    input [1 : 0]                   AWBURST_in_MD_CL2;
    input [1 : 0]                   AWLOCK_in_MD_CL2;
    input [3 : 0]                   AWCACHE_in_MD_CL2;
    input [2 : 0]                   AWPROT_in_MD_CL2;
    input                           AWVALID_in_MD_CL2;
    output                          AWREADY_out_MD_CL2;
    input [3 : 0]                   WID_in_MD_CL2;
    input [63 : 0]                  WDATA_in_MD_CL2;
    input [7 : 0]                   WSTRB_in_MD_CL2;
    input                           WLAST_in_MD_CL2;
    input                           WVALID_in_MD_CL2;
    output                          WREADY_out_MD_CL2;
    output [3 : 0]                  BID_out_MD_CL2;
    output [1 : 0]                  BRESP_out_MD_CL2;
    output                          BVALID_out_MD_CL2;
    input                           BREADY_in_MD_CL2;
    input [3 : 0]                   ARID_in_MD_CL2;
    input [31 : 0]                  ARADDR_in_MD_CL2;
    input [7 : 0]                   ARLEN_in_MD_CL2;
    input [2 : 0]                   ARSIZE_in_MD_CL2;
    input [1 : 0]                   ARBURST_in_MD_CL2;
    input [1 : 0]                   ARLOCK_in_MD_CL2;
    input [3 : 0]                   ARCACHE_in_MD_CL2;
    input [2 : 0]                   ARPROT_in_MD_CL2;
    input                           ARVALID_in_MD_CL2;
    output                          ARREADY_out_MD_CL2;
    output [3 : 0]                  RID_out_MD_CL2;
    output [63 : 0]                 RDATA_out_MD_CL2;
    output [1 : 0]                  RRESP_out_MD_CL2;
    output                          RLAST_out_MD_CL2;
    output                          RVALID_out_MD_CL2;
    input                           RREADY_in_MD_CL2;
    input [`COUNTERWD - 1 : 0]      init_div_MD_CL2;
    input [3 : 0]                   AWID_in_MI_CL2;
    input [31 : 0]                  AWADDR_in_MI_CL2;
    input [7 : 0]                   AWLEN_in_MI_CL2;
    input [2 : 0]                   AWSIZE_in_MI_CL2;
    input [1 : 0]                   AWBURST_in_MI_CL2;
    input [1 : 0]                   AWLOCK_in_MI_CL2;
    input [3 : 0]                   AWCACHE_in_MI_CL2;
    input [2 : 0]                   AWPROT_in_MI_CL2;
    input                           AWVALID_in_MI_CL2;
    output                          AWREADY_out_MI_CL2;
    input [3 : 0]                   WID_in_MI_CL2;
    input [63 : 0]                  WDATA_in_MI_CL2;
    input [7 : 0]                   WSTRB_in_MI_CL2;
    input                           WLAST_in_MI_CL2;
    input                           WVALID_in_MI_CL2;
    output                          WREADY_out_MI_CL2;
    output [3 : 0]                  BID_out_MI_CL2;
    output [1 : 0]                  BRESP_out_MI_CL2;
    output                          BVALID_out_MI_CL2;
    input                           BREADY_in_MI_CL2;
    input [3 : 0]                   ARID_in_MI_CL2;
    input [31 : 0]                  ARADDR_in_MI_CL2;
    input [7 : 0]                   ARLEN_in_MI_CL2;
    input [2 : 0]                   ARSIZE_in_MI_CL2;
    input [1 : 0]                   ARBURST_in_MI_CL2;
    input [1 : 0]                   ARLOCK_in_MI_CL2;
    input [3 : 0]                   ARCACHE_in_MI_CL2;
    input [2 : 0]                   ARPROT_in_MI_CL2;
    input                           ARVALID_in_MI_CL2;
    output                          ARREADY_out_MI_CL2;
    output [3 : 0]                  RID_out_MI_CL2;
    output [63 : 0]                 RDATA_out_MI_CL2;
    output [1 : 0]                  RRESP_out_MI_CL2;
    output                          RLAST_out_MI_CL2;
    output                          RVALID_out_MI_CL2;
    input                           RREADY_in_MI_CL2;
    input [`COUNTERWD - 1 : 0]      init_div_MI_CL2;
    output [3 : 0]                  AWID_out_SD_CL2;
    output [31 : 0]                 AWADDR_out_SD_CL2;
    output [7 : 0]                  AWLEN_out_SD_CL2;
    output [2 : 0]                  AWSIZE_out_SD_CL2;
    output [1 : 0]                  AWBURST_out_SD_CL2;
    output [1 : 0]                  AWLOCK_out_SD_CL2;
    output [3 : 0]                  AWCACHE_out_SD_CL2;
    output [2 : 0]                  AWPROT_out_SD_CL2;
    output                          AWVALID_out_SD_CL2;
    input                           AWREADY_in_SD_CL2;
    output [3 : 0]                  WID_out_SD_CL2;
    output [63 : 0]                 WDATA_out_SD_CL2;
    output [7 : 0]                  WSTRB_out_SD_CL2;
    output                          WLAST_out_SD_CL2;
    output                          WVALID_out_SD_CL2;
    input                           WREADY_in_SD_CL2;
    input [3 : 0]                   BID_in_SD_CL2;
    input [1 : 0]                   BRESP_in_SD_CL2;
    input                           BVALID_in_SD_CL2;
    output                          BREADY_out_SD_CL2;
    output [3 : 0]                  ARID_out_SD_CL2;
    output [31 : 0]                 ARADDR_out_SD_CL2;
    output [7 : 0]                  ARLEN_out_SD_CL2;
    output [2 : 0]                  ARSIZE_out_SD_CL2;
    output [1 : 0]                  ARBURST_out_SD_CL2;
    output [1 : 0]                  ARLOCK_out_SD_CL2;
    output [3 : 0]                  ARCACHE_out_SD_CL2;
    output [2 : 0]                  ARPROT_out_SD_CL2;
    output                          ARVALID_out_SD_CL2;
    input                           ARREADY_in_SD_CL2;
    input [3 : 0]                   RID_in_SD_CL2;
    input [63 : 0]                  RDATA_in_SD_CL2;
    input [1 : 0]                   RRESP_in_SD_CL2;
    input                           RLAST_in_SD_CL2;
    input                           RVALID_in_SD_CL2;
    output                          RREADY_out_SD_CL2;
    input [`COUNTERWD - 1 : 0]      target_div_SD_CL2;
    input [3 : 0]                   AWID_in_MD_CL3;
    input [31 : 0]                  AWADDR_in_MD_CL3;
    input [7 : 0]                   AWLEN_in_MD_CL3;
    input [2 : 0]                   AWSIZE_in_MD_CL3;
    input [1 : 0]                   AWBURST_in_MD_CL3;
    input [1 : 0]                   AWLOCK_in_MD_CL3;
    input [3 : 0]                   AWCACHE_in_MD_CL3;
    input [2 : 0]                   AWPROT_in_MD_CL3;
    input                           AWVALID_in_MD_CL3;
    output                          AWREADY_out_MD_CL3;
    input [3 : 0]                   WID_in_MD_CL3;
    input [63 : 0]                  WDATA_in_MD_CL3;
    input [7 : 0]                   WSTRB_in_MD_CL3;
    input                           WLAST_in_MD_CL3;
    input                           WVALID_in_MD_CL3;
    output                          WREADY_out_MD_CL3;
    output [3 : 0]                  BID_out_MD_CL3;
    output [1 : 0]                  BRESP_out_MD_CL3;
    output                          BVALID_out_MD_CL3;
    input                           BREADY_in_MD_CL3;
    input [3 : 0]                   ARID_in_MD_CL3;
    input [31 : 0]                  ARADDR_in_MD_CL3;
    input [7 : 0]                   ARLEN_in_MD_CL3;
    input [2 : 0]                   ARSIZE_in_MD_CL3;
    input [1 : 0]                   ARBURST_in_MD_CL3;
    input [1 : 0]                   ARLOCK_in_MD_CL3;
    input [3 : 0]                   ARCACHE_in_MD_CL3;
    input [2 : 0]                   ARPROT_in_MD_CL3;
    input                           ARVALID_in_MD_CL3;
    output                          ARREADY_out_MD_CL3;
    output [3 : 0]                  RID_out_MD_CL3;
    output [63 : 0]                 RDATA_out_MD_CL3;
    output [1 : 0]                  RRESP_out_MD_CL3;
    output                          RLAST_out_MD_CL3;
    output                          RVALID_out_MD_CL3;
    input                           RREADY_in_MD_CL3;
    input [`COUNTERWD - 1 : 0]      init_div_MD_CL3;
    input [3 : 0]                   AWID_in_MI_CL3;
    input [31 : 0]                  AWADDR_in_MI_CL3;
    input [7 : 0]                   AWLEN_in_MI_CL3;
    input [2 : 0]                   AWSIZE_in_MI_CL3;
    input [1 : 0]                   AWBURST_in_MI_CL3;
    input [1 : 0]                   AWLOCK_in_MI_CL3;
    input [3 : 0]                   AWCACHE_in_MI_CL3;
    input [2 : 0]                   AWPROT_in_MI_CL3;
    input                           AWVALID_in_MI_CL3;
    output                          AWREADY_out_MI_CL3;
    input [3 : 0]                   WID_in_MI_CL3;
    input [63 : 0]                  WDATA_in_MI_CL3;
    input [7 : 0]                   WSTRB_in_MI_CL3;
    input                           WLAST_in_MI_CL3;
    input                           WVALID_in_MI_CL3;
    output                          WREADY_out_MI_CL3;
    output [3 : 0]                  BID_out_MI_CL3;
    output [1 : 0]                  BRESP_out_MI_CL3;
    output                          BVALID_out_MI_CL3;
    input                           BREADY_in_MI_CL3;
    input [3 : 0]                   ARID_in_MI_CL3;
    input [31 : 0]                  ARADDR_in_MI_CL3;
    input [7 : 0]                   ARLEN_in_MI_CL3;
    input [2 : 0]                   ARSIZE_in_MI_CL3;
    input [1 : 0]                   ARBURST_in_MI_CL3;
    input [1 : 0]                   ARLOCK_in_MI_CL3;
    input [3 : 0]                   ARCACHE_in_MI_CL3;
    input [2 : 0]                   ARPROT_in_MI_CL3;
    input                           ARVALID_in_MI_CL3;
    output                          ARREADY_out_MI_CL3;
    output [3 : 0]                  RID_out_MI_CL3;
    output [63 : 0]                 RDATA_out_MI_CL3;
    output [1 : 0]                  RRESP_out_MI_CL3;
    output                          RLAST_out_MI_CL3;
    output                          RVALID_out_MI_CL3;
    input                           RREADY_in_MI_CL3;
    input [`COUNTERWD - 1 : 0]      init_div_MI_CL3;
    output [3 : 0]                  AWID_out_SD_CL3;
    output [31 : 0]                 AWADDR_out_SD_CL3;
    output [7 : 0]                  AWLEN_out_SD_CL3;
    output [2 : 0]                  AWSIZE_out_SD_CL3;
    output [1 : 0]                  AWBURST_out_SD_CL3;
    output [1 : 0]                  AWLOCK_out_SD_CL3;
    output [3 : 0]                  AWCACHE_out_SD_CL3;
    output [2 : 0]                  AWPROT_out_SD_CL3;
    output                          AWVALID_out_SD_CL3;
    input                           AWREADY_in_SD_CL3;
    output [3 : 0]                  WID_out_SD_CL3;
    output [63 : 0]                 WDATA_out_SD_CL3;
    output [7 : 0]                  WSTRB_out_SD_CL3;
    output                          WLAST_out_SD_CL3;
    output                          WVALID_out_SD_CL3;
    input                           WREADY_in_SD_CL3;
    input [3 : 0]                   BID_in_SD_CL3;
    input [1 : 0]                   BRESP_in_SD_CL3;
    input                           BVALID_in_SD_CL3;
    output                          BREADY_out_SD_CL3;
    output [3 : 0]                  ARID_out_SD_CL3;
    output [31 : 0]                 ARADDR_out_SD_CL3;
    output [7 : 0]                  ARLEN_out_SD_CL3;
    output [2 : 0]                  ARSIZE_out_SD_CL3;
    output [1 : 0]                  ARBURST_out_SD_CL3;
    output [1 : 0]                  ARLOCK_out_SD_CL3;
    output [3 : 0]                  ARCACHE_out_SD_CL3;
    output [2 : 0]                  ARPROT_out_SD_CL3;
    output                          ARVALID_out_SD_CL3;
    input                           ARREADY_in_SD_CL3;
    input [3 : 0]                   RID_in_SD_CL3;
    input [63 : 0]                  RDATA_in_SD_CL3;
    input [1 : 0]                   RRESP_in_SD_CL3;
    input                           RLAST_in_SD_CL3;
    input                           RVALID_in_SD_CL3;
    output                          RREADY_out_SD_CL3;
    input [`COUNTERWD - 1 : 0]      target_div_SD_CL3;
    output [3 : 0]                  AWID_out_L2_MEM;
    output [31 : 0]                 AWADDR_out_L2_MEM;
    output [7 : 0]                  AWLEN_out_L2_MEM;
    output [2 : 0]                  AWSIZE_out_L2_MEM;
    output [1 : 0]                  AWBURST_out_L2_MEM;
    output [1 : 0]                  AWLOCK_out_L2_MEM;
    output [3 : 0]                  AWCACHE_out_L2_MEM;
    output [2 : 0]                  AWPROT_out_L2_MEM;
    output                          AWVALID_out_L2_MEM;
    input                           AWREADY_in_L2_MEM;
    output [3 : 0]                  WID_out_L2_MEM;
    output [63 : 0]                 WDATA_out_L2_MEM;
    output [7 : 0]                  WSTRB_out_L2_MEM;
    output                          WLAST_out_L2_MEM;
    output                          WVALID_out_L2_MEM;
    input                           WREADY_in_L2_MEM;
    input [3 : 0]                   BID_in_L2_MEM;
    input [1 : 0]                   BRESP_in_L2_MEM;
    input                           BVALID_in_L2_MEM;
    output                          BREADY_out_L2_MEM;
    output [3 : 0]                  ARID_out_L2_MEM;
    output [31 : 0]                 ARADDR_out_L2_MEM;
    output [7 : 0]                  ARLEN_out_L2_MEM;
    output [2 : 0]                  ARSIZE_out_L2_MEM;
    output [1 : 0]                  ARBURST_out_L2_MEM;
    output [1 : 0]                  ARLOCK_out_L2_MEM;
    output [3 : 0]                  ARCACHE_out_L2_MEM;
    output [2 : 0]                  ARPROT_out_L2_MEM;
    output                          ARVALID_out_L2_MEM;
    input                           ARREADY_in_L2_MEM;
    input [3 : 0]                   RID_in_L2_MEM;
    input [63 : 0]                  RDATA_in_L2_MEM;
    input [1 : 0]                   RRESP_in_L2_MEM;
    input                           RLAST_in_L2_MEM;
    input                           RVALID_in_L2_MEM;
    output                          RREADY_out_L2_MEM;
    input [`COUNTERWD - 1 : 0]      target_div_L2_MEM;
    input [3 : 0]                   AWID_in_EXT;
    input [31 : 0]                  AWADDR_in_EXT;
    input [7 : 0]                   AWLEN_in_EXT;
    input [2 : 0]                   AWSIZE_in_EXT;
    input [1 : 0]                   AWBURST_in_EXT;
    input [1 : 0]                   AWLOCK_in_EXT;
    input [3 : 0]                   AWCACHE_in_EXT;
    input [2 : 0]                   AWPROT_in_EXT;
    input                           AWVALID_in_EXT;
    output                          AWREADY_out_EXT;
    input [3 : 0]                   WID_in_EXT;
    input [63 : 0]                  WDATA_in_EXT;
    input [7 : 0]                   WSTRB_in_EXT;
    input                           WLAST_in_EXT;
    input                           WVALID_in_EXT;
    output                          WREADY_out_EXT;
    output [3 : 0]                  BID_out_EXT;
    output [1 : 0]                  BRESP_out_EXT;
    output                          BVALID_out_EXT;
    input                           BREADY_in_EXT;
    input [3 : 0]                   ARID_in_EXT;
    input [31 : 0]                  ARADDR_in_EXT;
    input [7 : 0]                   ARLEN_in_EXT;
    input [2 : 0]                   ARSIZE_in_EXT;
    input [1 : 0]                   ARBURST_in_EXT;
    input [1 : 0]                   ARLOCK_in_EXT;
    input [3 : 0]                   ARCACHE_in_EXT;
    input [2 : 0]                   ARPROT_in_EXT;
    input                           ARVALID_in_EXT;
    output                          ARREADY_out_EXT;
    output [3 : 0]                  RID_out_EXT;
    output [63 : 0]                 RDATA_out_EXT;
    output [1 : 0]                  RRESP_out_EXT;
    output                          RLAST_out_EXT;
    output                          RVALID_out_EXT;
    input                           RREADY_in_EXT;
    input [`COUNTERWD - 1 : 0]      init_div_EXT;


    // Wires across switches
    wire signal_BWDAUX1_318767514_0;
    wire signal_BWDAUX2_318767514_0;
    wire signal_BWDAUX3_318767514_0;
    wire [79 : 0] signal_FLIT_318767514_0;
    wire signal_VALID_318767514_0;
    wire signal_FWDAUX1_318767514_0;
    wire signal_BWDAUX1_318767515_0;
    wire signal_BWDAUX2_318767515_0;
    wire signal_BWDAUX3_318767515_0;
    wire [79 : 0] signal_FLIT_318767515_0;
    wire signal_VALID_318767515_0;
    wire signal_FWDAUX1_318767515_0;
    wire signal_BWDAUX1_318767516_0;
    wire signal_BWDAUX2_318767516_0;
    wire signal_BWDAUX3_318767516_0;
    wire [79 : 0] signal_FLIT_318767516_0;
    wire signal_VALID_318767516_0;
    wire signal_FWDAUX1_318767516_0;
    wire signal_BWDAUX1_318767517_0;
    wire signal_BWDAUX2_318767517_0;
    wire signal_BWDAUX3_318767517_0;
    wire [79 : 0] signal_FLIT_318767517_0;
    wire signal_VALID_318767517_0;
    wire signal_FWDAUX1_318767517_0;
    wire signal_BWDAUX1_318767518_0;
    wire signal_BWDAUX2_318767518_0;
    wire signal_BWDAUX3_318767518_0;
    wire [79 : 0] signal_FLIT_318767518_0;
    wire signal_VALID_318767518_0;
    wire signal_FWDAUX1_318767518_0;
    wire signal_BWDAUX1_318767519_0;
    wire signal_BWDAUX2_318767519_0;
    wire signal_BWDAUX3_318767519_0;
    wire [79 : 0] signal_FLIT_318767519_0;
    wire signal_VALID_318767519_0;
    wire signal_FWDAUX1_318767519_0;
    wire signal_BWDAUX1_318767520_0;
    wire signal_BWDAUX2_318767520_0;
    wire signal_BWDAUX3_318767520_0;
    wire [79 : 0] signal_FLIT_318767520_0;
    wire signal_VALID_318767520_0;
    wire signal_FWDAUX1_318767520_0;
    wire signal_BWDAUX1_318767521_0;
    wire signal_BWDAUX2_318767521_0;
    wire signal_BWDAUX3_318767521_0;
    wire [79 : 0] signal_FLIT_318767521_0;
    wire signal_VALID_318767521_0;
    wire signal_FWDAUX1_318767521_0;
    wire signal_BWDAUX1_318767522_0;
    wire signal_BWDAUX2_318767522_0;
    wire signal_BWDAUX3_318767522_0;
    wire [79 : 0] signal_FLIT_318767522_0;
    wire signal_VALID_318767522_0;
    wire signal_FWDAUX1_318767522_0;
    wire signal_BWDAUX1_318767523_0;
    wire signal_BWDAUX2_318767523_0;
    wire signal_BWDAUX3_318767523_0;
    wire [79 : 0] signal_FLIT_318767523_0;
    wire signal_VALID_318767523_0;
    wire signal_FWDAUX1_318767523_0;
    wire signal_BWDAUX1_318767524_0;
    wire signal_BWDAUX2_318767524_0;
    wire signal_BWDAUX3_318767524_0;
    wire [79 : 0] signal_FLIT_318767524_0;
    wire signal_VALID_318767524_0;
    wire signal_FWDAUX1_318767524_0;
    wire signal_BWDAUX1_318767525_0;
    wire signal_BWDAUX2_318767525_0;
    wire signal_BWDAUX3_318767525_0;
    wire [79 : 0] signal_FLIT_318767525_0;
    wire signal_VALID_318767525_0;
    wire signal_FWDAUX1_318767525_0;
    wire signal_BWDAUX1_318767526_0;
    wire signal_BWDAUX2_318767526_0;
    wire signal_BWDAUX3_318767526_0;
    wire [79 : 0] signal_FLIT_318767526_0;
    wire signal_VALID_318767526_0;
    wire signal_FWDAUX1_318767526_0;
    wire signal_BWDAUX1_318767527_0;
    wire signal_BWDAUX2_318767527_0;
    wire signal_BWDAUX3_318767527_0;
    wire [79 : 0] signal_FLIT_318767527_0;
    wire signal_VALID_318767527_0;
    wire signal_FWDAUX1_318767527_0;
    wire signal_BWDAUX1_318767528_0;
    wire signal_BWDAUX2_318767528_0;
    wire signal_BWDAUX3_318767528_0;
    wire [79 : 0] signal_FLIT_318767528_0;
    wire signal_VALID_318767528_0;
    wire signal_FWDAUX1_318767528_0;
    wire signal_BWDAUX1_318767529_0;
    wire signal_BWDAUX2_318767529_0;
    wire signal_BWDAUX3_318767529_0;
    wire [79 : 0] signal_FLIT_318767529_0;
    wire signal_VALID_318767529_0;
    wire signal_FWDAUX1_318767529_0;
    wire signal_BWDAUX1_318767530_0;
    wire signal_BWDAUX2_318767530_0;
    wire signal_BWDAUX3_318767530_0;
    wire [79 : 0] signal_FLIT_318767530_0;
    wire signal_VALID_318767530_0;
    wire signal_FWDAUX1_318767530_0;
    wire signal_BWDAUX1_318767531_0;
    wire signal_BWDAUX2_318767531_0;
    wire signal_BWDAUX3_318767531_0;
    wire [79 : 0] signal_FLIT_318767531_0;
    wire signal_VALID_318767531_0;
    wire signal_FWDAUX1_318767531_0;
    wire signal_BWDAUX1_318767532_0;
    wire signal_BWDAUX2_318767532_0;
    wire signal_BWDAUX3_318767532_0;
    wire [79 : 0] signal_FLIT_318767532_0;
    wire signal_VALID_318767532_0;
    wire signal_FWDAUX1_318767532_0;
    wire signal_BWDAUX1_318767533_0;
    wire signal_BWDAUX2_318767533_0;
    wire signal_BWDAUX3_318767533_0;
    wire [79 : 0] signal_FLIT_318767533_0;
    wire signal_VALID_318767533_0;
    wire signal_FWDAUX1_318767533_0;
    wire signal_BWDAUX1_318767534_0;
    wire signal_BWDAUX2_318767534_0;
    wire signal_BWDAUX3_318767534_0;
    wire [79 : 0] signal_FLIT_318767534_0;
    wire signal_VALID_318767534_0;
    wire signal_FWDAUX1_318767534_0;
    wire signal_BWDAUX1_318767535_0;
    wire signal_BWDAUX2_318767535_0;
    wire signal_BWDAUX3_318767535_0;
    wire [79 : 0] signal_FLIT_318767535_0;
    wire signal_VALID_318767535_0;
    wire signal_FWDAUX1_318767535_0;
    wire signal_BWDAUX1_318767536_0;
    wire signal_BWDAUX2_318767536_0;
    wire signal_BWDAUX3_318767536_0;
    wire [79 : 0] signal_FLIT_318767536_0;
    wire signal_VALID_318767536_0;
    wire signal_FWDAUX1_318767536_0;
    wire signal_BWDAUX1_318767537_0;
    wire signal_BWDAUX2_318767537_0;
    wire signal_BWDAUX3_318767537_0;
    wire [79 : 0] signal_FLIT_318767537_0;
    wire signal_VALID_318767537_0;
    wire signal_FWDAUX1_318767537_0;
    wire signal_BWDAUX1_318767538_0;
    wire signal_BWDAUX2_318767538_0;
    wire signal_BWDAUX3_318767538_0;
    wire [79 : 0] signal_FLIT_318767538_0;
    wire signal_VALID_318767538_0;
    wire signal_FWDAUX1_318767538_0;
    wire signal_BWDAUX1_318767539_0;
    wire signal_BWDAUX2_318767539_0;
    wire signal_BWDAUX3_318767539_0;
    wire [79 : 0] signal_FLIT_318767539_0;
    wire signal_VALID_318767539_0;
    wire signal_FWDAUX1_318767539_0;
    wire signal_BWDAUX1_318767540_0;
    wire signal_BWDAUX2_318767540_0;
    wire signal_BWDAUX3_318767540_0;
    wire [79 : 0] signal_FLIT_318767540_0;
    wire signal_VALID_318767540_0;
    wire signal_FWDAUX1_318767540_0;
    wire signal_BWDAUX1_318767541_0;
    wire signal_BWDAUX2_318767541_0;
    wire signal_BWDAUX3_318767541_0;
    wire [79 : 0] signal_FLIT_318767541_0;
    wire signal_VALID_318767541_0;
    wire signal_FWDAUX1_318767541_0;
    wire signal_BWDAUX1_318767542_0;
    wire signal_BWDAUX2_318767542_0;
    wire signal_BWDAUX3_318767542_0;
    wire [79 : 0] signal_FLIT_318767542_0;
    wire signal_VALID_318767542_0;
    wire signal_FWDAUX1_318767542_0;
    wire signal_BWDAUX1_318767543_0;
    wire signal_BWDAUX2_318767543_0;
    wire signal_BWDAUX3_318767543_0;
    wire [79 : 0] signal_FLIT_318767543_0;
    wire signal_VALID_318767543_0;
    wire signal_FWDAUX1_318767543_0;
    wire signal_BWDAUX1_318767544_0;
    wire signal_BWDAUX2_318767544_0;
    wire signal_BWDAUX3_318767544_0;
    wire [79 : 0] signal_FLIT_318767544_0;
    wire signal_VALID_318767544_0;
    wire signal_FWDAUX1_318767544_0;
    wire signal_BWDAUX1_318767545_0;
    wire signal_BWDAUX2_318767545_0;
    wire signal_BWDAUX3_318767545_0;
    wire [79 : 0] signal_FLIT_318767545_0;
    wire signal_VALID_318767545_0;
    wire signal_FWDAUX1_318767545_0;
    
    ni_initiator_67109005_CLUSTER_0 ni_initiator_67109005(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MD_CL0), .rst(rst), .FLIT_in(signal_FLIT_318767538_0), .VALID_in(signal_VALID_318767538_0), .FWDAUX1_in(signal_FWDAUX1_318767538_0), .BWDAUX1_out(signal_BWDAUX1_318767538_0), .BWDAUX2_out(signal_BWDAUX2_318767538_0), .BWDAUX3_out(signal_BWDAUX3_318767538_0), .FLIT_out(signal_FLIT_318767528_0), .VALID_out(signal_VALID_318767528_0), .FWDAUX1_out(signal_FWDAUX1_318767528_0), .BWDAUX1_in(signal_BWDAUX1_318767528_0), .BWDAUX2_in(signal_BWDAUX2_318767528_0), .BWDAUX3_in(signal_BWDAUX3_318767528_0), .AWID(AWID_in_MD_CL0), .AWADDR(AWADDR_in_MD_CL0), .AWLEN(AWLEN_in_MD_CL0), .AWSIZE(AWSIZE_in_MD_CL0), .AWBURST(AWBURST_in_MD_CL0), .AWLOCK(AWLOCK_in_MD_CL0), .AWCACHE(AWCACHE_in_MD_CL0), .AWPROT(AWPROT_in_MD_CL0), .AWVALID(AWVALID_in_MD_CL0), .AWREADY(AWREADY_out_MD_CL0), .WID(WID_in_MD_CL0), .WDATA(WDATA_in_MD_CL0), .WSTRB(WSTRB_in_MD_CL0), .WLAST(WLAST_in_MD_CL0), .WVALID(WVALID_in_MD_CL0), .WREADY(WREADY_out_MD_CL0), .ARID(ARID_in_MD_CL0), .ARADDR(ARADDR_in_MD_CL0), .ARLEN(ARLEN_in_MD_CL0), .ARSIZE(ARSIZE_in_MD_CL0), .ARBURST(ARBURST_in_MD_CL0), .ARLOCK(ARLOCK_in_MD_CL0), .ARCACHE(ARCACHE_in_MD_CL0), .ARPROT(ARPROT_in_MD_CL0), .ARVALID(ARVALID_in_MD_CL0), .ARREADY(ARREADY_out_MD_CL0), .RID(RID_out_MD_CL0), .RDATA(RDATA_out_MD_CL0), .RRESP(RRESP_out_MD_CL0), .RLAST(RLAST_out_MD_CL0), .RVALID(RVALID_out_MD_CL0), .RREADY(RREADY_in_MD_CL0), .BID(BID_out_MD_CL0), .BRESP(BRESP_out_MD_CL0), .BVALID(BVALID_out_MD_CL0), .BREADY(BREADY_in_MD_CL0));

    ni_target_67109006_CLUSTER_0 ni_target_67109006(.core_clk(clk), .noc_clk(clk), .Clock_div(target_div_SD_CL0), .rst(rst), .FLIT_in(signal_FLIT_318767532_0), .VALID_in(signal_VALID_318767532_0), .FWDAUX1_in(signal_FWDAUX1_318767532_0), .BWDAUX1_out(signal_BWDAUX1_318767532_0), .BWDAUX2_out(signal_BWDAUX2_318767532_0), .BWDAUX3_out(signal_BWDAUX3_318767532_0), .FLIT_out(signal_FLIT_318767535_0), .VALID_out(signal_VALID_318767535_0), .FWDAUX1_out(signal_FWDAUX1_318767535_0), .BWDAUX1_in(signal_BWDAUX1_318767535_0), .BWDAUX2_in(signal_BWDAUX2_318767535_0), .BWDAUX3_in(signal_BWDAUX3_318767535_0), .AWID(AWID_out_SD_CL0), .AWADDR(AWADDR_out_SD_CL0), .AWLEN(AWLEN_out_SD_CL0), .AWSIZE(AWSIZE_out_SD_CL0), .AWBURST(AWBURST_out_SD_CL0), .AWLOCK(AWLOCK_out_SD_CL0), .AWCACHE(AWCACHE_out_SD_CL0), .AWPROT(AWPROT_out_SD_CL0), .AWVALID(AWVALID_out_SD_CL0), .AWREADY(AWREADY_in_SD_CL0), .WID(WID_out_SD_CL0), .WDATA(WDATA_out_SD_CL0), .WSTRB(WSTRB_out_SD_CL0), .WLAST(WLAST_out_SD_CL0), .WVALID(WVALID_out_SD_CL0), .WREADY(WREADY_in_SD_CL0), .ARID(ARID_out_SD_CL0), .ARADDR(ARADDR_out_SD_CL0), .ARLEN(ARLEN_out_SD_CL0), .ARSIZE(ARSIZE_out_SD_CL0), .ARBURST(ARBURST_out_SD_CL0), .ARLOCK(ARLOCK_out_SD_CL0), .ARCACHE(ARCACHE_out_SD_CL0), .ARPROT(ARPROT_out_SD_CL0), .ARVALID(ARVALID_out_SD_CL0), .ARREADY(ARREADY_in_SD_CL0), .RID(RID_in_SD_CL0), .RDATA(RDATA_in_SD_CL0), .RRESP(RRESP_in_SD_CL0), .RLAST(RLAST_in_SD_CL0), .RVALID(RVALID_in_SD_CL0), .RREADY(RREADY_out_SD_CL0), .BID(BID_in_SD_CL0), .BRESP(BRESP_in_SD_CL0), .BVALID(BVALID_in_SD_CL0), .BREADY(BREADY_out_SD_CL0));

    ni_initiator_67109007_CLUSTER_0 ni_initiator_67109007(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MI_CL0), .rst(rst), .FLIT_in(signal_FLIT_318767523_0), .VALID_in(signal_VALID_318767523_0), .FWDAUX1_in(signal_FWDAUX1_318767523_0), .BWDAUX1_out(signal_BWDAUX1_318767523_0), .BWDAUX2_out(signal_BWDAUX2_318767523_0), .BWDAUX3_out(signal_BWDAUX3_318767523_0), .FLIT_out(signal_FLIT_318767514_0), .VALID_out(signal_VALID_318767514_0), .FWDAUX1_out(signal_FWDAUX1_318767514_0), .BWDAUX1_in(signal_BWDAUX1_318767514_0), .BWDAUX2_in(signal_BWDAUX2_318767514_0), .BWDAUX3_in(signal_BWDAUX3_318767514_0), .AWID(AWID_in_MI_CL0), .AWADDR(AWADDR_in_MI_CL0), .AWLEN(AWLEN_in_MI_CL0), .AWSIZE(AWSIZE_in_MI_CL0), .AWBURST(AWBURST_in_MI_CL0), .AWLOCK(AWLOCK_in_MI_CL0), .AWCACHE(AWCACHE_in_MI_CL0), .AWPROT(AWPROT_in_MI_CL0), .AWVALID(AWVALID_in_MI_CL0), .AWREADY(AWREADY_out_MI_CL0), .WID(WID_in_MI_CL0), .WDATA(WDATA_in_MI_CL0), .WSTRB(WSTRB_in_MI_CL0), .WLAST(WLAST_in_MI_CL0), .WVALID(WVALID_in_MI_CL0), .WREADY(WREADY_out_MI_CL0), .ARID(ARID_in_MI_CL0), .ARADDR(ARADDR_in_MI_CL0), .ARLEN(ARLEN_in_MI_CL0), .ARSIZE(ARSIZE_in_MI_CL0), .ARBURST(ARBURST_in_MI_CL0), .ARLOCK(ARLOCK_in_MI_CL0), .ARCACHE(ARCACHE_in_MI_CL0), .ARPROT(ARPROT_in_MI_CL0), .ARVALID(ARVALID_in_MI_CL0), .ARREADY(ARREADY_out_MI_CL0), .RID(RID_out_MI_CL0), .RDATA(RDATA_out_MI_CL0), .RRESP(RRESP_out_MI_CL0), .RLAST(RLAST_out_MI_CL0), .RVALID(RVALID_out_MI_CL0), .RREADY(RREADY_in_MI_CL0), .BID(BID_out_MI_CL0), .BRESP(BRESP_out_MI_CL0), .BVALID(BVALID_out_MI_CL0), .BREADY(BREADY_in_MI_CL0));

    ni_initiator_67109008_CLUSTER_1 ni_initiator_67109008(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MD_CL1), .rst(rst), .FLIT_in(signal_FLIT_318767539_0), .VALID_in(signal_VALID_318767539_0), .FWDAUX1_in(signal_FWDAUX1_318767539_0), .BWDAUX1_out(signal_BWDAUX1_318767539_0), .BWDAUX2_out(signal_BWDAUX2_318767539_0), .BWDAUX3_out(signal_BWDAUX3_318767539_0), .FLIT_out(signal_FLIT_318767529_0), .VALID_out(signal_VALID_318767529_0), .FWDAUX1_out(signal_FWDAUX1_318767529_0), .BWDAUX1_in(signal_BWDAUX1_318767529_0), .BWDAUX2_in(signal_BWDAUX2_318767529_0), .BWDAUX3_in(signal_BWDAUX3_318767529_0), .AWID(AWID_in_MD_CL1), .AWADDR(AWADDR_in_MD_CL1), .AWLEN(AWLEN_in_MD_CL1), .AWSIZE(AWSIZE_in_MD_CL1), .AWBURST(AWBURST_in_MD_CL1), .AWLOCK(AWLOCK_in_MD_CL1), .AWCACHE(AWCACHE_in_MD_CL1), .AWPROT(AWPROT_in_MD_CL1), .AWVALID(AWVALID_in_MD_CL1), .AWREADY(AWREADY_out_MD_CL1), .WID(WID_in_MD_CL1), .WDATA(WDATA_in_MD_CL1), .WSTRB(WSTRB_in_MD_CL1), .WLAST(WLAST_in_MD_CL1), .WVALID(WVALID_in_MD_CL1), .WREADY(WREADY_out_MD_CL1), .ARID(ARID_in_MD_CL1), .ARADDR(ARADDR_in_MD_CL1), .ARLEN(ARLEN_in_MD_CL1), .ARSIZE(ARSIZE_in_MD_CL1), .ARBURST(ARBURST_in_MD_CL1), .ARLOCK(ARLOCK_in_MD_CL1), .ARCACHE(ARCACHE_in_MD_CL1), .ARPROT(ARPROT_in_MD_CL1), .ARVALID(ARVALID_in_MD_CL1), .ARREADY(ARREADY_out_MD_CL1), .RID(RID_out_MD_CL1), .RDATA(RDATA_out_MD_CL1), .RRESP(RRESP_out_MD_CL1), .RLAST(RLAST_out_MD_CL1), .RVALID(RVALID_out_MD_CL1), .RREADY(RREADY_in_MD_CL1), .BID(BID_out_MD_CL1), .BRESP(BRESP_out_MD_CL1), .BVALID(BVALID_out_MD_CL1), .BREADY(BREADY_in_MD_CL1));

    ni_initiator_67109009_CLUSTER_1 ni_initiator_67109009(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MI_CL1), .rst(rst), .FLIT_in(signal_FLIT_318767524_0), .VALID_in(signal_VALID_318767524_0), .FWDAUX1_in(signal_FWDAUX1_318767524_0), .BWDAUX1_out(signal_BWDAUX1_318767524_0), .BWDAUX2_out(signal_BWDAUX2_318767524_0), .BWDAUX3_out(signal_BWDAUX3_318767524_0), .FLIT_out(signal_FLIT_318767515_0), .VALID_out(signal_VALID_318767515_0), .FWDAUX1_out(signal_FWDAUX1_318767515_0), .BWDAUX1_in(signal_BWDAUX1_318767515_0), .BWDAUX2_in(signal_BWDAUX2_318767515_0), .BWDAUX3_in(signal_BWDAUX3_318767515_0), .AWID(AWID_in_MI_CL1), .AWADDR(AWADDR_in_MI_CL1), .AWLEN(AWLEN_in_MI_CL1), .AWSIZE(AWSIZE_in_MI_CL1), .AWBURST(AWBURST_in_MI_CL1), .AWLOCK(AWLOCK_in_MI_CL1), .AWCACHE(AWCACHE_in_MI_CL1), .AWPROT(AWPROT_in_MI_CL1), .AWVALID(AWVALID_in_MI_CL1), .AWREADY(AWREADY_out_MI_CL1), .WID(WID_in_MI_CL1), .WDATA(WDATA_in_MI_CL1), .WSTRB(WSTRB_in_MI_CL1), .WLAST(WLAST_in_MI_CL1), .WVALID(WVALID_in_MI_CL1), .WREADY(WREADY_out_MI_CL1), .ARID(ARID_in_MI_CL1), .ARADDR(ARADDR_in_MI_CL1), .ARLEN(ARLEN_in_MI_CL1), .ARSIZE(ARSIZE_in_MI_CL1), .ARBURST(ARBURST_in_MI_CL1), .ARLOCK(ARLOCK_in_MI_CL1), .ARCACHE(ARCACHE_in_MI_CL1), .ARPROT(ARPROT_in_MI_CL1), .ARVALID(ARVALID_in_MI_CL1), .ARREADY(ARREADY_out_MI_CL1), .RID(RID_out_MI_CL1), .RDATA(RDATA_out_MI_CL1), .RRESP(RRESP_out_MI_CL1), .RLAST(RLAST_out_MI_CL1), .RVALID(RVALID_out_MI_CL1), .RREADY(RREADY_in_MI_CL1), .BID(BID_out_MI_CL1), .BRESP(BRESP_out_MI_CL1), .BVALID(BVALID_out_MI_CL1), .BREADY(BREADY_in_MI_CL1));

    ni_target_67109010_CLUSTER_1 ni_target_67109010(.core_clk(clk), .noc_clk(clk), .Clock_div(target_div_SD_CL1), .rst(rst), .FLIT_in(signal_FLIT_318767533_0), .VALID_in(signal_VALID_318767533_0), .FWDAUX1_in(signal_FWDAUX1_318767533_0), .BWDAUX1_out(signal_BWDAUX1_318767533_0), .BWDAUX2_out(signal_BWDAUX2_318767533_0), .BWDAUX3_out(signal_BWDAUX3_318767533_0), .FLIT_out(signal_FLIT_318767536_0), .VALID_out(signal_VALID_318767536_0), .FWDAUX1_out(signal_FWDAUX1_318767536_0), .BWDAUX1_in(signal_BWDAUX1_318767536_0), .BWDAUX2_in(signal_BWDAUX2_318767536_0), .BWDAUX3_in(signal_BWDAUX3_318767536_0), .AWID(AWID_out_SD_CL1), .AWADDR(AWADDR_out_SD_CL1), .AWLEN(AWLEN_out_SD_CL1), .AWSIZE(AWSIZE_out_SD_CL1), .AWBURST(AWBURST_out_SD_CL1), .AWLOCK(AWLOCK_out_SD_CL1), .AWCACHE(AWCACHE_out_SD_CL1), .AWPROT(AWPROT_out_SD_CL1), .AWVALID(AWVALID_out_SD_CL1), .AWREADY(AWREADY_in_SD_CL1), .WID(WID_out_SD_CL1), .WDATA(WDATA_out_SD_CL1), .WSTRB(WSTRB_out_SD_CL1), .WLAST(WLAST_out_SD_CL1), .WVALID(WVALID_out_SD_CL1), .WREADY(WREADY_in_SD_CL1), .ARID(ARID_out_SD_CL1), .ARADDR(ARADDR_out_SD_CL1), .ARLEN(ARLEN_out_SD_CL1), .ARSIZE(ARSIZE_out_SD_CL1), .ARBURST(ARBURST_out_SD_CL1), .ARLOCK(ARLOCK_out_SD_CL1), .ARCACHE(ARCACHE_out_SD_CL1), .ARPROT(ARPROT_out_SD_CL1), .ARVALID(ARVALID_out_SD_CL1), .ARREADY(ARREADY_in_SD_CL1), .RID(RID_in_SD_CL1), .RDATA(RDATA_in_SD_CL1), .RRESP(RRESP_in_SD_CL1), .RLAST(RLAST_in_SD_CL1), .RVALID(RVALID_in_SD_CL1), .RREADY(RREADY_out_SD_CL1), .BID(BID_in_SD_CL1), .BRESP(BRESP_in_SD_CL1), .BVALID(BVALID_in_SD_CL1), .BREADY(BREADY_out_SD_CL1));

    ni_initiator_67109011_CLUSTER_2 ni_initiator_67109011(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MD_CL2), .rst(rst), .FLIT_in(signal_FLIT_318767540_0), .VALID_in(signal_VALID_318767540_0), .FWDAUX1_in(signal_FWDAUX1_318767540_0), .BWDAUX1_out(signal_BWDAUX1_318767540_0), .BWDAUX2_out(signal_BWDAUX2_318767540_0), .BWDAUX3_out(signal_BWDAUX3_318767540_0), .FLIT_out(signal_FLIT_318767530_0), .VALID_out(signal_VALID_318767530_0), .FWDAUX1_out(signal_FWDAUX1_318767530_0), .BWDAUX1_in(signal_BWDAUX1_318767530_0), .BWDAUX2_in(signal_BWDAUX2_318767530_0), .BWDAUX3_in(signal_BWDAUX3_318767530_0), .AWID(AWID_in_MD_CL2), .AWADDR(AWADDR_in_MD_CL2), .AWLEN(AWLEN_in_MD_CL2), .AWSIZE(AWSIZE_in_MD_CL2), .AWBURST(AWBURST_in_MD_CL2), .AWLOCK(AWLOCK_in_MD_CL2), .AWCACHE(AWCACHE_in_MD_CL2), .AWPROT(AWPROT_in_MD_CL2), .AWVALID(AWVALID_in_MD_CL2), .AWREADY(AWREADY_out_MD_CL2), .WID(WID_in_MD_CL2), .WDATA(WDATA_in_MD_CL2), .WSTRB(WSTRB_in_MD_CL2), .WLAST(WLAST_in_MD_CL2), .WVALID(WVALID_in_MD_CL2), .WREADY(WREADY_out_MD_CL2), .ARID(ARID_in_MD_CL2), .ARADDR(ARADDR_in_MD_CL2), .ARLEN(ARLEN_in_MD_CL2), .ARSIZE(ARSIZE_in_MD_CL2), .ARBURST(ARBURST_in_MD_CL2), .ARLOCK(ARLOCK_in_MD_CL2), .ARCACHE(ARCACHE_in_MD_CL2), .ARPROT(ARPROT_in_MD_CL2), .ARVALID(ARVALID_in_MD_CL2), .ARREADY(ARREADY_out_MD_CL2), .RID(RID_out_MD_CL2), .RDATA(RDATA_out_MD_CL2), .RRESP(RRESP_out_MD_CL2), .RLAST(RLAST_out_MD_CL2), .RVALID(RVALID_out_MD_CL2), .RREADY(RREADY_in_MD_CL2), .BID(BID_out_MD_CL2), .BRESP(BRESP_out_MD_CL2), .BVALID(BVALID_out_MD_CL2), .BREADY(BREADY_in_MD_CL2));

    ni_initiator_67109012_CLUSTER_2 ni_initiator_67109012(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MI_CL2), .rst(rst), .FLIT_in(signal_FLIT_318767525_0), .VALID_in(signal_VALID_318767525_0), .FWDAUX1_in(signal_FWDAUX1_318767525_0), .BWDAUX1_out(signal_BWDAUX1_318767525_0), .BWDAUX2_out(signal_BWDAUX2_318767525_0), .BWDAUX3_out(signal_BWDAUX3_318767525_0), .FLIT_out(signal_FLIT_318767516_0), .VALID_out(signal_VALID_318767516_0), .FWDAUX1_out(signal_FWDAUX1_318767516_0), .BWDAUX1_in(signal_BWDAUX1_318767516_0), .BWDAUX2_in(signal_BWDAUX2_318767516_0), .BWDAUX3_in(signal_BWDAUX3_318767516_0), .AWID(AWID_in_MI_CL2), .AWADDR(AWADDR_in_MI_CL2), .AWLEN(AWLEN_in_MI_CL2), .AWSIZE(AWSIZE_in_MI_CL2), .AWBURST(AWBURST_in_MI_CL2), .AWLOCK(AWLOCK_in_MI_CL2), .AWCACHE(AWCACHE_in_MI_CL2), .AWPROT(AWPROT_in_MI_CL2), .AWVALID(AWVALID_in_MI_CL2), .AWREADY(AWREADY_out_MI_CL2), .WID(WID_in_MI_CL2), .WDATA(WDATA_in_MI_CL2), .WSTRB(WSTRB_in_MI_CL2), .WLAST(WLAST_in_MI_CL2), .WVALID(WVALID_in_MI_CL2), .WREADY(WREADY_out_MI_CL2), .ARID(ARID_in_MI_CL2), .ARADDR(ARADDR_in_MI_CL2), .ARLEN(ARLEN_in_MI_CL2), .ARSIZE(ARSIZE_in_MI_CL2), .ARBURST(ARBURST_in_MI_CL2), .ARLOCK(ARLOCK_in_MI_CL2), .ARCACHE(ARCACHE_in_MI_CL2), .ARPROT(ARPROT_in_MI_CL2), .ARVALID(ARVALID_in_MI_CL2), .ARREADY(ARREADY_out_MI_CL2), .RID(RID_out_MI_CL2), .RDATA(RDATA_out_MI_CL2), .RRESP(RRESP_out_MI_CL2), .RLAST(RLAST_out_MI_CL2), .RVALID(RVALID_out_MI_CL2), .RREADY(RREADY_in_MI_CL2), .BID(BID_out_MI_CL2), .BRESP(BRESP_out_MI_CL2), .BVALID(BVALID_out_MI_CL2), .BREADY(BREADY_in_MI_CL2));

    ni_target_67109013_CLUSTER_2 ni_target_67109013(.core_clk(clk), .noc_clk(clk), .Clock_div(target_div_SD_CL2), .rst(rst), .FLIT_in(signal_FLIT_318767519_0), .VALID_in(signal_VALID_318767519_0), .FWDAUX1_in(signal_FWDAUX1_318767519_0), .BWDAUX1_out(signal_BWDAUX1_318767519_0), .BWDAUX2_out(signal_BWDAUX2_318767519_0), .BWDAUX3_out(signal_BWDAUX3_318767519_0), .FLIT_out(signal_FLIT_318767521_0), .VALID_out(signal_VALID_318767521_0), .FWDAUX1_out(signal_FWDAUX1_318767521_0), .BWDAUX1_in(signal_BWDAUX1_318767521_0), .BWDAUX2_in(signal_BWDAUX2_318767521_0), .BWDAUX3_in(signal_BWDAUX3_318767521_0), .AWID(AWID_out_SD_CL2), .AWADDR(AWADDR_out_SD_CL2), .AWLEN(AWLEN_out_SD_CL2), .AWSIZE(AWSIZE_out_SD_CL2), .AWBURST(AWBURST_out_SD_CL2), .AWLOCK(AWLOCK_out_SD_CL2), .AWCACHE(AWCACHE_out_SD_CL2), .AWPROT(AWPROT_out_SD_CL2), .AWVALID(AWVALID_out_SD_CL2), .AWREADY(AWREADY_in_SD_CL2), .WID(WID_out_SD_CL2), .WDATA(WDATA_out_SD_CL2), .WSTRB(WSTRB_out_SD_CL2), .WLAST(WLAST_out_SD_CL2), .WVALID(WVALID_out_SD_CL2), .WREADY(WREADY_in_SD_CL2), .ARID(ARID_out_SD_CL2), .ARADDR(ARADDR_out_SD_CL2), .ARLEN(ARLEN_out_SD_CL2), .ARSIZE(ARSIZE_out_SD_CL2), .ARBURST(ARBURST_out_SD_CL2), .ARLOCK(ARLOCK_out_SD_CL2), .ARCACHE(ARCACHE_out_SD_CL2), .ARPROT(ARPROT_out_SD_CL2), .ARVALID(ARVALID_out_SD_CL2), .ARREADY(ARREADY_in_SD_CL2), .RID(RID_in_SD_CL2), .RDATA(RDATA_in_SD_CL2), .RRESP(RRESP_in_SD_CL2), .RLAST(RLAST_in_SD_CL2), .RVALID(RVALID_in_SD_CL2), .RREADY(RREADY_out_SD_CL2), .BID(BID_in_SD_CL2), .BRESP(BRESP_in_SD_CL2), .BVALID(BVALID_in_SD_CL2), .BREADY(BREADY_out_SD_CL2));

    ni_initiator_67109014_CLUSTER_3 ni_initiator_67109014(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MD_CL3), .rst(rst), .FLIT_in(signal_FLIT_318767526_0), .VALID_in(signal_VALID_318767526_0), .FWDAUX1_in(signal_FWDAUX1_318767526_0), .BWDAUX1_out(signal_BWDAUX1_318767526_0), .BWDAUX2_out(signal_BWDAUX2_318767526_0), .BWDAUX3_out(signal_BWDAUX3_318767526_0), .FLIT_out(signal_FLIT_318767517_0), .VALID_out(signal_VALID_318767517_0), .FWDAUX1_out(signal_FWDAUX1_318767517_0), .BWDAUX1_in(signal_BWDAUX1_318767517_0), .BWDAUX2_in(signal_BWDAUX2_318767517_0), .BWDAUX3_in(signal_BWDAUX3_318767517_0), .AWID(AWID_in_MD_CL3), .AWADDR(AWADDR_in_MD_CL3), .AWLEN(AWLEN_in_MD_CL3), .AWSIZE(AWSIZE_in_MD_CL3), .AWBURST(AWBURST_in_MD_CL3), .AWLOCK(AWLOCK_in_MD_CL3), .AWCACHE(AWCACHE_in_MD_CL3), .AWPROT(AWPROT_in_MD_CL3), .AWVALID(AWVALID_in_MD_CL3), .AWREADY(AWREADY_out_MD_CL3), .WID(WID_in_MD_CL3), .WDATA(WDATA_in_MD_CL3), .WSTRB(WSTRB_in_MD_CL3), .WLAST(WLAST_in_MD_CL3), .WVALID(WVALID_in_MD_CL3), .WREADY(WREADY_out_MD_CL3), .ARID(ARID_in_MD_CL3), .ARADDR(ARADDR_in_MD_CL3), .ARLEN(ARLEN_in_MD_CL3), .ARSIZE(ARSIZE_in_MD_CL3), .ARBURST(ARBURST_in_MD_CL3), .ARLOCK(ARLOCK_in_MD_CL3), .ARCACHE(ARCACHE_in_MD_CL3), .ARPROT(ARPROT_in_MD_CL3), .ARVALID(ARVALID_in_MD_CL3), .ARREADY(ARREADY_out_MD_CL3), .RID(RID_out_MD_CL3), .RDATA(RDATA_out_MD_CL3), .RRESP(RRESP_out_MD_CL3), .RLAST(RLAST_out_MD_CL3), .RVALID(RVALID_out_MD_CL3), .RREADY(RREADY_in_MD_CL3), .BID(BID_out_MD_CL3), .BRESP(BRESP_out_MD_CL3), .BVALID(BVALID_out_MD_CL3), .BREADY(BREADY_in_MD_CL3));

    ni_initiator_67109015_CLUSTER_3 ni_initiator_67109015(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_MI_CL3), .rst(rst), .FLIT_in(signal_FLIT_318767527_0), .VALID_in(signal_VALID_318767527_0), .FWDAUX1_in(signal_FWDAUX1_318767527_0), .BWDAUX1_out(signal_BWDAUX1_318767527_0), .BWDAUX2_out(signal_BWDAUX2_318767527_0), .BWDAUX3_out(signal_BWDAUX3_318767527_0), .FLIT_out(signal_FLIT_318767518_0), .VALID_out(signal_VALID_318767518_0), .FWDAUX1_out(signal_FWDAUX1_318767518_0), .BWDAUX1_in(signal_BWDAUX1_318767518_0), .BWDAUX2_in(signal_BWDAUX2_318767518_0), .BWDAUX3_in(signal_BWDAUX3_318767518_0), .AWID(AWID_in_MI_CL3), .AWADDR(AWADDR_in_MI_CL3), .AWLEN(AWLEN_in_MI_CL3), .AWSIZE(AWSIZE_in_MI_CL3), .AWBURST(AWBURST_in_MI_CL3), .AWLOCK(AWLOCK_in_MI_CL3), .AWCACHE(AWCACHE_in_MI_CL3), .AWPROT(AWPROT_in_MI_CL3), .AWVALID(AWVALID_in_MI_CL3), .AWREADY(AWREADY_out_MI_CL3), .WID(WID_in_MI_CL3), .WDATA(WDATA_in_MI_CL3), .WSTRB(WSTRB_in_MI_CL3), .WLAST(WLAST_in_MI_CL3), .WVALID(WVALID_in_MI_CL3), .WREADY(WREADY_out_MI_CL3), .ARID(ARID_in_MI_CL3), .ARADDR(ARADDR_in_MI_CL3), .ARLEN(ARLEN_in_MI_CL3), .ARSIZE(ARSIZE_in_MI_CL3), .ARBURST(ARBURST_in_MI_CL3), .ARLOCK(ARLOCK_in_MI_CL3), .ARCACHE(ARCACHE_in_MI_CL3), .ARPROT(ARPROT_in_MI_CL3), .ARVALID(ARVALID_in_MI_CL3), .ARREADY(ARREADY_out_MI_CL3), .RID(RID_out_MI_CL3), .RDATA(RDATA_out_MI_CL3), .RRESP(RRESP_out_MI_CL3), .RLAST(RLAST_out_MI_CL3), .RVALID(RVALID_out_MI_CL3), .RREADY(RREADY_in_MI_CL3), .BID(BID_out_MI_CL3), .BRESP(BRESP_out_MI_CL3), .BVALID(BVALID_out_MI_CL3), .BREADY(BREADY_in_MI_CL3));

    ni_target_67109016_CLUSTER_3 ni_target_67109016(.core_clk(clk), .noc_clk(clk), .Clock_div(target_div_SD_CL3), .rst(rst), .FLIT_in(signal_FLIT_318767534_0), .VALID_in(signal_VALID_318767534_0), .FWDAUX1_in(signal_FWDAUX1_318767534_0), .BWDAUX1_out(signal_BWDAUX1_318767534_0), .BWDAUX2_out(signal_BWDAUX2_318767534_0), .BWDAUX3_out(signal_BWDAUX3_318767534_0), .FLIT_out(signal_FLIT_318767537_0), .VALID_out(signal_VALID_318767537_0), .FWDAUX1_out(signal_FWDAUX1_318767537_0), .BWDAUX1_in(signal_BWDAUX1_318767537_0), .BWDAUX2_in(signal_BWDAUX2_318767537_0), .BWDAUX3_in(signal_BWDAUX3_318767537_0), .AWID(AWID_out_SD_CL3), .AWADDR(AWADDR_out_SD_CL3), .AWLEN(AWLEN_out_SD_CL3), .AWSIZE(AWSIZE_out_SD_CL3), .AWBURST(AWBURST_out_SD_CL3), .AWLOCK(AWLOCK_out_SD_CL3), .AWCACHE(AWCACHE_out_SD_CL3), .AWPROT(AWPROT_out_SD_CL3), .AWVALID(AWVALID_out_SD_CL3), .AWREADY(AWREADY_in_SD_CL3), .WID(WID_out_SD_CL3), .WDATA(WDATA_out_SD_CL3), .WSTRB(WSTRB_out_SD_CL3), .WLAST(WLAST_out_SD_CL3), .WVALID(WVALID_out_SD_CL3), .WREADY(WREADY_in_SD_CL3), .ARID(ARID_out_SD_CL3), .ARADDR(ARADDR_out_SD_CL3), .ARLEN(ARLEN_out_SD_CL3), .ARSIZE(ARSIZE_out_SD_CL3), .ARBURST(ARBURST_out_SD_CL3), .ARLOCK(ARLOCK_out_SD_CL3), .ARCACHE(ARCACHE_out_SD_CL3), .ARPROT(ARPROT_out_SD_CL3), .ARVALID(ARVALID_out_SD_CL3), .ARREADY(ARREADY_in_SD_CL3), .RID(RID_in_SD_CL3), .RDATA(RDATA_in_SD_CL3), .RRESP(RRESP_in_SD_CL3), .RLAST(RLAST_in_SD_CL3), .RVALID(RVALID_in_SD_CL3), .RREADY(RREADY_out_SD_CL3), .BID(BID_in_SD_CL3), .BRESP(BRESP_in_SD_CL3), .BVALID(BVALID_in_SD_CL3), .BREADY(BREADY_out_SD_CL3));

    ni_target_67109017_L2_MEM ni_target_67109017(.core_clk(clk), .noc_clk(clk), .Clock_div(target_div_L2_MEM), .rst(rst), .FLIT_in(signal_FLIT_318767520_0), .VALID_in(signal_VALID_318767520_0), .FWDAUX1_in(signal_FWDAUX1_318767520_0), .BWDAUX1_out(signal_BWDAUX1_318767520_0), .BWDAUX2_out(signal_BWDAUX2_318767520_0), .BWDAUX3_out(signal_BWDAUX3_318767520_0), .FLIT_out(signal_FLIT_318767522_0), .VALID_out(signal_VALID_318767522_0), .FWDAUX1_out(signal_FWDAUX1_318767522_0), .BWDAUX1_in(signal_BWDAUX1_318767522_0), .BWDAUX2_in(signal_BWDAUX2_318767522_0), .BWDAUX3_in(signal_BWDAUX3_318767522_0), .AWID(AWID_out_L2_MEM), .AWADDR(AWADDR_out_L2_MEM), .AWLEN(AWLEN_out_L2_MEM), .AWSIZE(AWSIZE_out_L2_MEM), .AWBURST(AWBURST_out_L2_MEM), .AWLOCK(AWLOCK_out_L2_MEM), .AWCACHE(AWCACHE_out_L2_MEM), .AWPROT(AWPROT_out_L2_MEM), .AWVALID(AWVALID_out_L2_MEM), .AWREADY(AWREADY_in_L2_MEM), .WID(WID_out_L2_MEM), .WDATA(WDATA_out_L2_MEM), .WSTRB(WSTRB_out_L2_MEM), .WLAST(WLAST_out_L2_MEM), .WVALID(WVALID_out_L2_MEM), .WREADY(WREADY_in_L2_MEM), .ARID(ARID_out_L2_MEM), .ARADDR(ARADDR_out_L2_MEM), .ARLEN(ARLEN_out_L2_MEM), .ARSIZE(ARSIZE_out_L2_MEM), .ARBURST(ARBURST_out_L2_MEM), .ARLOCK(ARLOCK_out_L2_MEM), .ARCACHE(ARCACHE_out_L2_MEM), .ARPROT(ARPROT_out_L2_MEM), .ARVALID(ARVALID_out_L2_MEM), .ARREADY(ARREADY_in_L2_MEM), .RID(RID_in_L2_MEM), .RDATA(RDATA_in_L2_MEM), .RRESP(RRESP_in_L2_MEM), .RLAST(RLAST_in_L2_MEM), .RVALID(RVALID_in_L2_MEM), .RREADY(RREADY_out_L2_MEM), .BID(BID_in_L2_MEM), .BRESP(BRESP_in_L2_MEM), .BVALID(BVALID_in_L2_MEM), .BREADY(BREADY_out_L2_MEM));

    ni_initiator_67109018_SOC_MASTER ni_initiator_67109018(.core_clk(clk), .noc_clk(clk), .Clock_div(init_div_EXT), .rst(rst), .FLIT_in(signal_FLIT_318767541_0), .VALID_in(signal_VALID_318767541_0), .FWDAUX1_in(signal_FWDAUX1_318767541_0), .BWDAUX1_out(signal_BWDAUX1_318767541_0), .BWDAUX2_out(signal_BWDAUX2_318767541_0), .BWDAUX3_out(signal_BWDAUX3_318767541_0), .FLIT_out(signal_FLIT_318767531_0), .VALID_out(signal_VALID_318767531_0), .FWDAUX1_out(signal_FWDAUX1_318767531_0), .BWDAUX1_in(signal_BWDAUX1_318767531_0), .BWDAUX2_in(signal_BWDAUX2_318767531_0), .BWDAUX3_in(signal_BWDAUX3_318767531_0), .AWID(AWID_in_EXT), .AWADDR(AWADDR_in_EXT), .AWLEN(AWLEN_in_EXT), .AWSIZE(AWSIZE_in_EXT), .AWBURST(AWBURST_in_EXT), .AWLOCK(AWLOCK_in_EXT), .AWCACHE(AWCACHE_in_EXT), .AWPROT(AWPROT_in_EXT), .AWVALID(AWVALID_in_EXT), .AWREADY(AWREADY_out_EXT), .WID(WID_in_EXT), .WDATA(WDATA_in_EXT), .WSTRB(WSTRB_in_EXT), .WLAST(WLAST_in_EXT), .WVALID(WVALID_in_EXT), .WREADY(WREADY_out_EXT), .ARID(ARID_in_EXT), .ARADDR(ARADDR_in_EXT), .ARLEN(ARLEN_in_EXT), .ARSIZE(ARSIZE_in_EXT), .ARBURST(ARBURST_in_EXT), .ARLOCK(ARLOCK_in_EXT), .ARCACHE(ARCACHE_in_EXT), .ARPROT(ARPROT_in_EXT), .ARVALID(ARVALID_in_EXT), .ARREADY(ARREADY_out_EXT), .RID(RID_out_EXT), .RDATA(RDATA_out_EXT), .RRESP(RRESP_out_EXT), .RLAST(RLAST_out_EXT), .RVALID(RVALID_out_EXT), .RREADY(RREADY_in_EXT), .BID(BID_out_EXT), .BRESP(BRESP_out_EXT), .BVALID(BVALID_out_EXT), .BREADY(BREADY_in_EXT));

    switch_16777291 sw_16777291(.clk(clk), .rst(rst), .FLIT_in_0(signal_FLIT_318767514_0), .VALID_in_0(signal_VALID_318767514_0), .FWDAUX1_in_0(signal_FWDAUX1_318767514_0), .BWDAUX1_out_0(signal_BWDAUX1_318767514_0), .BWDAUX2_out_0(signal_BWDAUX2_318767514_0), .BWDAUX3_out_0(signal_BWDAUX3_318767514_0), .FLIT_in_1(signal_FLIT_318767515_0), .VALID_in_1(signal_VALID_318767515_0), .FWDAUX1_in_1(signal_FWDAUX1_318767515_0), .BWDAUX1_out_1(signal_BWDAUX1_318767515_0), .BWDAUX2_out_1(signal_BWDAUX2_318767515_0), .BWDAUX3_out_1(signal_BWDAUX3_318767515_0), .FLIT_in_2(signal_FLIT_318767516_0), .VALID_in_2(signal_VALID_318767516_0), .FWDAUX1_in_2(signal_FWDAUX1_318767516_0), .BWDAUX1_out_2(signal_BWDAUX1_318767516_0), .BWDAUX2_out_2(signal_BWDAUX2_318767516_0), .BWDAUX3_out_2(signal_BWDAUX3_318767516_0), .FLIT_in_3(signal_FLIT_318767517_0), .VALID_in_3(signal_VALID_318767517_0), .FWDAUX1_in_3(signal_FWDAUX1_318767517_0), .BWDAUX1_out_3(signal_BWDAUX1_318767517_0), .BWDAUX2_out_3(signal_BWDAUX2_318767517_0), .BWDAUX3_out_3(signal_BWDAUX3_318767517_0), .FLIT_in_4(signal_FLIT_318767518_0), .VALID_in_4(signal_VALID_318767518_0), .FWDAUX1_in_4(signal_FWDAUX1_318767518_0), .BWDAUX1_out_4(signal_BWDAUX1_318767518_0), .BWDAUX2_out_4(signal_BWDAUX2_318767518_0), .BWDAUX3_out_4(signal_BWDAUX3_318767518_0), .FLIT_in_5(signal_FLIT_318767542_0), .VALID_in_5(signal_VALID_318767542_0), .FWDAUX1_in_5(signal_FWDAUX1_318767542_0), .BWDAUX1_out_5(signal_BWDAUX1_318767542_0), .BWDAUX2_out_5(signal_BWDAUX2_318767542_0), .BWDAUX3_out_5(signal_BWDAUX3_318767542_0), .FLIT_out_0(signal_FLIT_318767519_0), .VALID_out_0(signal_VALID_318767519_0), .FWDAUX1_out_0(signal_FWDAUX1_318767519_0), .BWDAUX1_in_0(signal_BWDAUX1_318767519_0), .BWDAUX2_in_0(signal_BWDAUX2_318767519_0), .BWDAUX3_in_0(signal_BWDAUX3_318767519_0), .FLIT_out_1(signal_FLIT_318767520_0), .VALID_out_1(signal_VALID_318767520_0), .FWDAUX1_out_1(signal_FWDAUX1_318767520_0), .BWDAUX1_in_1(signal_BWDAUX1_318767520_0), .BWDAUX2_in_1(signal_BWDAUX2_318767520_0), .BWDAUX3_in_1(signal_BWDAUX3_318767520_0), .FLIT_out_2(signal_FLIT_318767543_0), .VALID_out_2(signal_VALID_318767543_0), .FWDAUX1_out_2(signal_FWDAUX1_318767543_0), .BWDAUX1_in_2(signal_BWDAUX1_318767543_0), .BWDAUX2_in_2(signal_BWDAUX2_318767543_0), .BWDAUX3_in_2(signal_BWDAUX3_318767543_0));
    
    switch_16777292 sw_16777292(.clk(clk), .rst(rst), .FLIT_in_0(signal_FLIT_318767521_0), .VALID_in_0(signal_VALID_318767521_0), .FWDAUX1_in_0(signal_FWDAUX1_318767521_0), .BWDAUX1_out_0(signal_BWDAUX1_318767521_0), .BWDAUX2_out_0(signal_BWDAUX2_318767521_0), .BWDAUX3_out_0(signal_BWDAUX3_318767521_0), .FLIT_in_1(signal_FLIT_318767522_0), .VALID_in_1(signal_VALID_318767522_0), .FWDAUX1_in_1(signal_FWDAUX1_318767522_0), .BWDAUX1_out_1(signal_BWDAUX1_318767522_0), .BWDAUX2_out_1(signal_BWDAUX2_318767522_0), .BWDAUX3_out_1(signal_BWDAUX3_318767522_0), .FLIT_in_2(signal_FLIT_318767545_0), .VALID_in_2(signal_VALID_318767545_0), .FWDAUX1_in_2(signal_FWDAUX1_318767545_0), .BWDAUX1_out_2(signal_BWDAUX1_318767545_0), .BWDAUX2_out_2(signal_BWDAUX2_318767545_0), .BWDAUX3_out_2(signal_BWDAUX3_318767545_0), .FLIT_out_0(signal_FLIT_318767523_0), .VALID_out_0(signal_VALID_318767523_0), .FWDAUX1_out_0(signal_FWDAUX1_318767523_0), .BWDAUX1_in_0(signal_BWDAUX1_318767523_0), .BWDAUX2_in_0(signal_BWDAUX2_318767523_0), .BWDAUX3_in_0(signal_BWDAUX3_318767523_0), .FLIT_out_1(signal_FLIT_318767524_0), .VALID_out_1(signal_VALID_318767524_0), .FWDAUX1_out_1(signal_FWDAUX1_318767524_0), .BWDAUX1_in_1(signal_BWDAUX1_318767524_0), .BWDAUX2_in_1(signal_BWDAUX2_318767524_0), .BWDAUX3_in_1(signal_BWDAUX3_318767524_0), .FLIT_out_2(signal_FLIT_318767525_0), .VALID_out_2(signal_VALID_318767525_0), .FWDAUX1_out_2(signal_FWDAUX1_318767525_0), .BWDAUX1_in_2(signal_BWDAUX1_318767525_0), .BWDAUX2_in_2(signal_BWDAUX2_318767525_0), .BWDAUX3_in_2(signal_BWDAUX3_318767525_0), .FLIT_out_3(signal_FLIT_318767526_0), .VALID_out_3(signal_VALID_318767526_0), .FWDAUX1_out_3(signal_FWDAUX1_318767526_0), .BWDAUX1_in_3(signal_BWDAUX1_318767526_0), .BWDAUX2_in_3(signal_BWDAUX2_318767526_0), .BWDAUX3_in_3(signal_BWDAUX3_318767526_0), .FLIT_out_4(signal_FLIT_318767527_0), .VALID_out_4(signal_VALID_318767527_0), .FWDAUX1_out_4(signal_FWDAUX1_318767527_0), .BWDAUX1_in_4(signal_BWDAUX1_318767527_0), .BWDAUX2_in_4(signal_BWDAUX2_318767527_0), .BWDAUX3_in_4(signal_BWDAUX3_318767527_0), .FLIT_out_5(signal_FLIT_318767544_0), .VALID_out_5(signal_VALID_318767544_0), .FWDAUX1_out_5(signal_FWDAUX1_318767544_0), .BWDAUX1_in_5(signal_BWDAUX1_318767544_0), .BWDAUX2_in_5(signal_BWDAUX2_318767544_0), .BWDAUX3_in_5(signal_BWDAUX3_318767544_0));
    
    switch_16777293 sw_16777293(.clk(clk), .rst(rst), .FLIT_in_0(signal_FLIT_318767528_0), .VALID_in_0(signal_VALID_318767528_0), .FWDAUX1_in_0(signal_FWDAUX1_318767528_0), .BWDAUX1_out_0(signal_BWDAUX1_318767528_0), .BWDAUX2_out_0(signal_BWDAUX2_318767528_0), .BWDAUX3_out_0(signal_BWDAUX3_318767528_0), .FLIT_in_1(signal_FLIT_318767529_0), .VALID_in_1(signal_VALID_318767529_0), .FWDAUX1_in_1(signal_FWDAUX1_318767529_0), .BWDAUX1_out_1(signal_BWDAUX1_318767529_0), .BWDAUX2_out_1(signal_BWDAUX2_318767529_0), .BWDAUX3_out_1(signal_BWDAUX3_318767529_0), .FLIT_in_2(signal_FLIT_318767530_0), .VALID_in_2(signal_VALID_318767530_0), .FWDAUX1_in_2(signal_FWDAUX1_318767530_0), .BWDAUX1_out_2(signal_BWDAUX1_318767530_0), .BWDAUX2_out_2(signal_BWDAUX2_318767530_0), .BWDAUX3_out_2(signal_BWDAUX3_318767530_0), .FLIT_in_3(signal_FLIT_318767531_0), .VALID_in_3(signal_VALID_318767531_0), .FWDAUX1_in_3(signal_FWDAUX1_318767531_0), .BWDAUX1_out_3(signal_BWDAUX1_318767531_0), .BWDAUX2_out_3(signal_BWDAUX2_318767531_0), .BWDAUX3_out_3(signal_BWDAUX3_318767531_0), .FLIT_in_4(signal_FLIT_318767543_0), .VALID_in_4(signal_VALID_318767543_0), .FWDAUX1_in_4(signal_FWDAUX1_318767543_0), .BWDAUX1_out_4(signal_BWDAUX1_318767543_0), .BWDAUX2_out_4(signal_BWDAUX2_318767543_0), .BWDAUX3_out_4(signal_BWDAUX3_318767543_0), .FLIT_out_0(signal_FLIT_318767532_0), .VALID_out_0(signal_VALID_318767532_0), .FWDAUX1_out_0(signal_FWDAUX1_318767532_0), .BWDAUX1_in_0(signal_BWDAUX1_318767532_0), .BWDAUX2_in_0(signal_BWDAUX2_318767532_0), .BWDAUX3_in_0(signal_BWDAUX3_318767532_0), .FLIT_out_1(signal_FLIT_318767533_0), .VALID_out_1(signal_VALID_318767533_0), .FWDAUX1_out_1(signal_FWDAUX1_318767533_0), .BWDAUX1_in_1(signal_BWDAUX1_318767533_0), .BWDAUX2_in_1(signal_BWDAUX2_318767533_0), .BWDAUX3_in_1(signal_BWDAUX3_318767533_0), .FLIT_out_2(signal_FLIT_318767534_0), .VALID_out_2(signal_VALID_318767534_0), .FWDAUX1_out_2(signal_FWDAUX1_318767534_0), .BWDAUX1_in_2(signal_BWDAUX1_318767534_0), .BWDAUX2_in_2(signal_BWDAUX2_318767534_0), .BWDAUX3_in_2(signal_BWDAUX3_318767534_0), .FLIT_out_3(signal_FLIT_318767542_0), .VALID_out_3(signal_VALID_318767542_0), .FWDAUX1_out_3(signal_FWDAUX1_318767542_0), .BWDAUX1_in_3(signal_BWDAUX1_318767542_0), .BWDAUX2_in_3(signal_BWDAUX2_318767542_0), .BWDAUX3_in_3(signal_BWDAUX3_318767542_0));
    
    switch_16777294 sw_16777294(.clk(clk), .rst(rst), .FLIT_in_0(signal_FLIT_318767535_0), .VALID_in_0(signal_VALID_318767535_0), .FWDAUX1_in_0(signal_FWDAUX1_318767535_0), .BWDAUX1_out_0(signal_BWDAUX1_318767535_0), .BWDAUX2_out_0(signal_BWDAUX2_318767535_0), .BWDAUX3_out_0(signal_BWDAUX3_318767535_0), .FLIT_in_1(signal_FLIT_318767536_0), .VALID_in_1(signal_VALID_318767536_0), .FWDAUX1_in_1(signal_FWDAUX1_318767536_0), .BWDAUX1_out_1(signal_BWDAUX1_318767536_0), .BWDAUX2_out_1(signal_BWDAUX2_318767536_0), .BWDAUX3_out_1(signal_BWDAUX3_318767536_0), .FLIT_in_2(signal_FLIT_318767537_0), .VALID_in_2(signal_VALID_318767537_0), .FWDAUX1_in_2(signal_FWDAUX1_318767537_0), .BWDAUX1_out_2(signal_BWDAUX1_318767537_0), .BWDAUX2_out_2(signal_BWDAUX2_318767537_0), .BWDAUX3_out_2(signal_BWDAUX3_318767537_0), .FLIT_in_3(signal_FLIT_318767544_0), .VALID_in_3(signal_VALID_318767544_0), .FWDAUX1_in_3(signal_FWDAUX1_318767544_0), .BWDAUX1_out_3(signal_BWDAUX1_318767544_0), .BWDAUX2_out_3(signal_BWDAUX2_318767544_0), .BWDAUX3_out_3(signal_BWDAUX3_318767544_0), .FLIT_out_0(signal_FLIT_318767538_0), .VALID_out_0(signal_VALID_318767538_0), .FWDAUX1_out_0(signal_FWDAUX1_318767538_0), .BWDAUX1_in_0(signal_BWDAUX1_318767538_0), .BWDAUX2_in_0(signal_BWDAUX2_318767538_0), .BWDAUX3_in_0(signal_BWDAUX3_318767538_0), .FLIT_out_1(signal_FLIT_318767539_0), .VALID_out_1(signal_VALID_318767539_0), .FWDAUX1_out_1(signal_FWDAUX1_318767539_0), .BWDAUX1_in_1(signal_BWDAUX1_318767539_0), .BWDAUX2_in_1(signal_BWDAUX2_318767539_0), .BWDAUX3_in_1(signal_BWDAUX3_318767539_0), .FLIT_out_2(signal_FLIT_318767540_0), .VALID_out_2(signal_VALID_318767540_0), .FWDAUX1_out_2(signal_FWDAUX1_318767540_0), .BWDAUX1_in_2(signal_BWDAUX1_318767540_0), .BWDAUX2_in_2(signal_BWDAUX2_318767540_0), .BWDAUX3_in_2(signal_BWDAUX3_318767540_0), .FLIT_out_3(signal_FLIT_318767541_0), .VALID_out_3(signal_VALID_318767541_0), .FWDAUX1_out_3(signal_FWDAUX1_318767541_0), .BWDAUX1_in_3(signal_BWDAUX1_318767541_0), .BWDAUX2_in_3(signal_BWDAUX2_318767541_0), .BWDAUX3_in_3(signal_BWDAUX3_318767541_0), .FLIT_out_4(signal_FLIT_318767545_0), .VALID_out_4(signal_VALID_318767545_0), .FWDAUX1_out_4(signal_FWDAUX1_318767545_0), .BWDAUX1_in_4(signal_BWDAUX1_318767545_0), .BWDAUX2_in_4(signal_BWDAUX2_318767545_0), .BWDAUX3_in_4(signal_BWDAUX3_318767545_0));
    
    
endmodule
