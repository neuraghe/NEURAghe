--!
--! @file fll_counter.vhd
--! @brief Frequency Locked Loop Counter 
--! 
--! This is the architecture model of the FLL counter.
--!
--! <B>
--! @n
--! This file is part of the Platform 2012 program,
--! a cooperation between STMicroelectronics and CEA.@n
--! Redistribution of this file to outside parties is
--! strictly prohibited without the written consent
--! of the module owner indicated below.@n
--! </B>
--! 
--! @par  Module owner: Pascal VIVET
--!       pascal.vivet@cea.fr
--! 
--! @par  Copyright (C) 2009 CEA
--! 
--! @par  Authors: Pascal VIVET
--! 
--! @par  Id: $Id: fll_counter.vhd 1 2014-01-15 16:11:08Z im219746 $
--! @par  Date: $Date: 2014-01-15 17:11:08 +0100 (Wed, 15 Jan 2014) $
--! @par  Revision: $Rev: 1 $
--!


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

LIBRARY common_cells_lib;
USE common_cells_lib.ALL;

ENTITY fll_counter IS
  PORT(
    clk_dco       : IN  STD_LOGIC;                    -- clk generated by the VCO/DCO
    rst_async_n   : IN  STD_LOGIC;                    -- hard reset
    test_mode     : IN  STD_LOGIC;                    -- test_mode from CVP-U
    clear         : IN  STD_LOGIC;                    -- counter clear (done by control unit when counter has been registered properly)
    sample_i      : IN  STD_LOGIC;                    -- sample input signal, set during NB cycles clk_ref
    sample_o      : OUT STD_LOGIC;                    -- sample output signal, resynchronized with clk_dco
    counter       : OUT STD_LOGIC_VECTOR(7 downto 0)  -- counter value, send back to control
    );
END fll_counter;

ARCHITECTURE rtl of fll_counter IS

  ----------------------------------------------------------------------
  -- Components declarations -------------------------------------------
  ----------------------------------------------------------------------

  COMPONENT reset_synchronizer IS
    GENERIC(
      SYNCHRONIZERS    : natural :=  5  -- Number of synchronizers 
    );
    PORT(
      clk        : IN  STD_LOGIC;
      rst_n      : IN  STD_LOGIC;
      test_mode  : IN  STD_LOGIC;

      rst_out_n  : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT clock_gating 
    PORT(
      clk_in      : IN  STD_LOGIC;
      enable      : IN  STD_LOGIC;
      test_mode   : IN  STD_LOGIC;
      clk_out     : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT clock_mux2 IS
    PORT(
      clk_in0     : IN  STD_LOGIC;
      clk_in1     : IN  STD_LOGIC;
      clk_select  : IN  STD_LOGIC;
  
      clk_out     : OUT STD_LOGIC
    );
  END COMPONENT;

  ----------------------------------------------------------------------
  -- Signals/contants declarations -------------------------------------
  ----------------------------------------------------------------------

  SIGNAL rst_resync_n    : STD_LOGIC;
  SIGNAL rst_or_clear_n  : STD_LOGIC;

  SIGNAL sample1, sample2, sample3, sample4 : STD_LOGIC;

  SIGNAL do_sample   : STD_LOGIC;

  SIGNAL counter_i   : STD_LOGIC_VECTOR(7 downto 0);
  SIGNAL counter_0   : STD_LOGIC;
  SIGNAL counter_0_s : STD_LOGIC;
  SIGNAL counter_1   : STD_LOGIC;
  SIGNAL counter_1_s : STD_LOGIC;

BEGIN

  --------------------------------------------------------------------------------
  -- reset resynchronization logic with clk_dco
  --------------------------------------------------------------------------------

  reset_resync_u: reset_synchronizer
    GENERIC MAP ( SYNCHRONIZERS => 2 )
    PORT MAP(
      clk        => clk_dco   ,
      rst_n      => rst_async_n,
      test_mode  => test_mode   ,
      rst_out_n  => rst_resync_n 
    );
  
  
  --------------------------------------------------------------------------------
  -- reset / clear signal of the counter :
  -- - use the clear signal from control unit : used as an asynchronous reset, active low during one 'clk' cycle
  --------------------------------------------------------------------------------

  rst_or_clear_n <= (not(clear) or test_mode) and rst_resync_n;
  
  
  --------------------------------------------------------------------------------
  -- sample signal resynchronization logic with clk_dco (4 stages sync due since at 4GHz - to be sure, who knows ...-)
  --------------------------------------------------------------------------------

  PROCESS (clk_dco, rst_resync_n)
  BEGIN
    IF (rst_resync_n = '0') THEN
      sample1 <= '0';
      sample2 <= '0';
      sample3 <= '0';
      sample4 <= '0';
    ELSIF clk_dco = '1' AND clk_dco'EVENT THEN
      sample1 <= sample_i;
      sample2 <= sample1;
      sample3 <= sample2;
      sample4 <= sample3;
    END IF;
  END PROCESS;


  --------------------------------------------------------------------------------
  -- asynchronous ripple adder : 1st stage
  --------------------------------------------------------------------------------
  
  -- the first stage clock is gated by the sample signal. Use proper clock gate element.
  u_do_sample_cg : clock_gating
    PORT MAP(
      clk_in      => clk_dco,
      enable      => sample4,
      test_mode   => test_mode,
      clk_out     => do_sample
    );
  
  PROCESS (do_sample, rst_or_clear_n)
  BEGIN
    IF (rst_or_clear_n = '0') THEN
      counter_0 <= '1';
    ELSIF do_sample = '1' AND do_sample'EVENT THEN  -- max freq ~ 4 GHz
        counter_0 <= not(counter_0);
    END IF;
  END PROCESS;

  counter_i(0) <= not(counter_0);  -- max freq ~ 2 GHz
  
  --------------------------------------------------------------------------------
  -- asynchronous ripple adder : 2nd stage
  --------------------------------------------------------------------------------
  
  clk_mux_for_test_counter_1_u : clock_mux2 
    PORT MAP(
      clk_in0     => counter_0,
      clk_in1     => clk_dco,
      clk_select  => test_mode,

      clk_out     => counter_0_s
    );
  
  PROCESS (counter_0_s, rst_or_clear_n)
  BEGIN
    IF (rst_or_clear_n = '0') THEN
      counter_1 <= '1';
    ELSIF counter_0_s = '1' AND counter_0_s'EVENT THEN  -- max freq ~ 2 GHz
      counter_1 <= not(counter_1);
    END IF;
  END PROCESS;

  counter_i(1) <= not(counter_1);  -- max freq ~ 1 GHz
  
  --------------------------------------------------------------------------------
  -- asynchronous ripple adder : standard 6 bit adder (7 downto 2)
  --------------------------------------------------------------------------------
  
  clk_mux_for_test_counters_u : clock_mux2 
    PORT MAP(
      clk_in0     => counter_1,
      clk_in1     => clk_dco,
      clk_select  => test_mode,

      clk_out     => counter_1_s
    );

  PROCESS (counter_1_s, rst_or_clear_n)
  BEGIN
    IF (rst_or_clear_n = '0') THEN
      counter_i(7 downto 2)   <= (others => '0');
    ELSIF counter_1_s = '1' AND counter_1_s'EVENT THEN    -- max freq ~ 1 GHz
      IF (counter_i(7 downto 2) /= "111111") THEN         -- avoid counter overflow
        counter_i(7 downto 2) <= UNSIGNED(counter_i(7 downto 2)) + 1;
      END IF;
    END IF;
  END PROCESS;


  --------------------------------------------------------------------------------
  -- output signals
  --------------------------------------------------------------------------------
  
  -- counter value
  counter <= counter_i;
  
  -- output count signal, resynchronized with clk_dco, in phase with the 'counter' output data.
  sample_o <= sample4;
  
END rtl;
