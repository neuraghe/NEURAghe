const logic [0:839][31:0] vector_out = {
32'h0cb20ccc,
32'h0ce60d00,
32'h0d1a0d34,
32'h0d4e0d68,
32'h0d820d9c,
32'h0db60dd0,
32'h0dea0e04,
32'h0e1e0e38,
32'h0e520e6c,
32'h0e860ea0,
32'h0eba0ed4,
32'h0eee0f08,
32'h0f220f3c,
32'h0f560f70,
32'h0f8a0fa4,
32'h0fbe0fd8,
32'h0ff2100c,
32'h10261040,
32'h105a1074,
32'h108e10a8,
32'h10c210dc,
32'h10f61110,
32'h112a1144,
32'h115e1178,
32'h119211ac,
32'h11c611e0,
32'h11fa1214,
32'h122e1248,
32'h1262127c,
32'h129612b0,
32'h132e1348,
32'h1362137c,
32'h139613b0,
32'h13ca13e4,
32'h13fe1418,
32'h1432144c,
32'h14661480,
32'h149a14b4,
32'h14ce14e8,
32'h1502151c,
32'h15361550,
32'h156a1584,
32'h159e15b8,
32'h15d215ec,
32'h16061620,
32'h163a1654,
32'h166e1688,
32'h16a216bc,
32'h16d616f0,
32'h170a1724,
32'h173e1758,
32'h1772178c,
32'h17a617c0,
32'h17da17f4,
32'h180e1828,
32'h1842185c,
32'h18761890,
32'h18aa18c4,
32'h18de18f8,
32'h1912192c,
32'h19aa19c4,
32'h19de19f8,
32'h1a121a2c,
32'h1a461a60,
32'h1a7a1a94,
32'h1aae1ac8,
32'h1ae21afc,
32'h1b161b30,
32'h1b4a1b64,
32'h1b7e1b98,
32'h1bb21bcc,
32'h1be61c00,
32'h1c1a1c34,
32'h1c4e1c68,
32'h1c821c9c,
32'h1cb61cd0,
32'h1cea1d04,
32'h1d1e1d38,
32'h1d521d6c,
32'h1d861da0,
32'h1dba1dd4,
32'h1dee1e08,
32'h1e221e3c,
32'h1e561e70,
32'h1e8a1ea4,
32'h1ebe1ed8,
32'h1ef21f0c,
32'h1f261f40,
32'h1f5a1f74,
32'h1f8e1fa8,
32'h20262040,
32'h205a2074,
32'h208e20a8,
32'h20c220dc,
32'h20f62110,
32'h212a2144,
32'h215e2178,
32'h219221ac,
32'h21c621e0,
32'h21fa2214,
32'h222e2248,
32'h2262227c,
32'h229622b0,
32'h22ca22e4,
32'h22fe2318,
32'h2332234c,
32'h23662380,
32'h239a23b4,
32'h23ce23e8,
32'h2402241c,
32'h24362450,
32'h246a2484,
32'h249e24b8,
32'h24d224ec,
32'h25062520,
32'h253a2554,
32'h256e2588,
32'h25a225bc,
32'h25d625f0,
32'h260a2624,
32'h26a226bc,
32'h26d626f0,
32'h270a2724,
32'h273e2758,
32'h2772278c,
32'h27a627c0,
32'h27da27f4,
32'h280e2828,
32'h2842285c,
32'h28762890,
32'h28aa28c4,
32'h28de28f8,
32'h2912292c,
32'h29462960,
32'h297a2994,
32'h29ae29c8,
32'h29e229fc,
32'h2a162a30,
32'h2a4a2a64,
32'h2a7e2a98,
32'h2ab22acc,
32'h2ae62b00,
32'h2b1a2b34,
32'h2b4e2b68,
32'h2b822b9c,
32'h2bb62bd0,
32'h2bea2c04,
32'h2c1e2c38,
32'h2c522c6c,
32'h2c862ca0,
32'h2d1e2d38,
32'h2d522d6c,
32'h2d862da0,
32'h2dba2dd4,
32'h2dee2e08,
32'h2e222e3c,
32'h2e562e70,
32'h2e8a2ea4,
32'h2ebe2ed8,
32'h2ef22f0c,
32'h2f262f40,
32'h2f5a2f74,
32'h2f8e2fa8,
32'h2fc22fdc,
32'h2ff63010,
32'h302a3044,
32'h305e3078,
32'h309230ac,
32'h30c630e0,
32'h30fa3114,
32'h312e3148,
32'h3162317c,
32'h319631b0,
32'h31ca31e4,
32'h31fe3218,
32'h3232324c,
32'h32663280,
32'h329a32b4,
32'h32ce32e8,
32'h3302331c,
32'h339a33b4,
32'h33ce33e8,
32'h3402341c,
32'h34363450,
32'h346a3484,
32'h349e34b8,
32'h34d234ec,
32'h35063520,
32'h353a3554,
32'h356e3588,
32'h35a235bc,
32'h35d635f0,
32'h360a3624,
32'h363e3658,
32'h3672368c,
32'h36a636c0,
32'h36da36f4,
32'h370e3728,
32'h3742375c,
32'h37763790,
32'h37aa37c4,
32'h37de37f8,
32'h3812382c,
32'h38463860,
32'h387a3894,
32'h38ae38c8,
32'h38e238fc,
32'h39163930,
32'h394a3964,
32'h397e3998,
32'h3a163a30,
32'h3a4a3a64,
32'h3a7e3a98,
32'h3ab23acc,
32'h3ae63b00,
32'h3b1a3b34,
32'h3b4e3b68,
32'h3b823b9c,
32'h3bb63bd0,
32'h3bea3c04,
32'h3c1e3c38,
32'h3c523c6c,
32'h3c863ca0,
32'h3cba3cd4,
32'h3cee3d08,
32'h3d223d3c,
32'h3d563d70,
32'h3d8a3da4,
32'h3dbe3dd8,
32'h3df23e0c,
32'h3e263e40,
32'h3e5a3e74,
32'h3e8e3ea8,
32'h3ec23edc,
32'h3ef63f10,
32'h3f2a3f44,
32'h3f5e3f78,
32'h3f923fac,
32'h3fc63fe0,
32'h3ffa4014,
32'h409240ac,
32'h40c640e0,
32'h40fa4114,
32'h412e4148,
32'h4162417c,
32'h419641b0,
32'h41ca41e4,
32'h41fe4218,
32'h4232424c,
32'h42664280,
32'h429a42b4,
32'h42ce42e8,
32'h4302431c,
32'h43364350,
32'h436a4384,
32'h439e43b8,
32'h43d243ec,
32'h44064420,
32'h443a4454,
32'h446e4488,
32'h44a244bc,
32'h44d644f0,
32'h450a4524,
32'h453e4558,
32'h4572458c,
32'h45a645c0,
32'h45da45f4,
32'h460e4628,
32'h4642465c,
32'h46764690,
32'h470e4728,
32'h4742475c,
32'h47764790,
32'h47aa47c4,
32'h47de47f8,
32'h4812482c,
32'h48464860,
32'h487a4894,
32'h48ae48c8,
32'h48e248fc,
32'h49164930,
32'h494a4964,
32'h497e4998,
32'h49b249cc,
32'h49e64a00,
32'h4a1a4a34,
32'h4a4e4a68,
32'h4a824a9c,
32'h4ab64ad0,
32'h4aea4b04,
32'h4b1e4b38,
32'h4b524b6c,
32'h4b864ba0,
32'h4bba4bd4,
32'h4bee4c08,
32'h4c224c3c,
32'h4c564c70,
32'h4c8a4ca4,
32'h4cbe4cd8,
32'h4cf24d0c,
32'h4d8a4da4,
32'h4dbe4dd8,
32'h4df24e0c,
32'h4e264e40,
32'h4e5a4e74,
32'h4e8e4ea8,
32'h4ec24edc,
32'h4ef64f10,
32'h4f2a4f44,
32'h4f5e4f78,
32'h4f924fac,
32'h4fc64fe0,
32'h4ffa5014,
32'h502e5048,
32'h5062507c,
32'h509650b0,
32'h50ca50e4,
32'h50fe5118,
32'h5132514c,
32'h51665180,
32'h519a51b4,
32'h51ce51e8,
32'h5202521c,
32'h52365250,
32'h526a5284,
32'h529e52b8,
32'h52d252ec,
32'h53065320,
32'h533a5354,
32'h536e5388,
32'h54065420,
32'h543a5454,
32'h546e5488,
32'h54a254bc,
32'h54d654f0,
32'h550a5524,
32'h553e5558,
32'h5572558c,
32'h55a655c0,
32'h55da55f4,
32'h560e5628,
32'h5642565c,
32'h56765690,
32'h56aa56c4,
32'h56de56f8,
32'h5712572c,
32'h57465760,
32'h577a5794,
32'h57ae57c8,
32'h57e257fc,
32'h58165830,
32'h584a5864,
32'h587e5898,
32'h58b258cc,
32'h58e65900,
32'h591a5934,
32'h594e5968,
32'h5982599c,
32'h59b659d0,
32'h59ea5a04,
32'h5a825a9c,
32'h5ab65ad0,
32'h5aea5b04,
32'h5b1e5b38,
32'h5b525b6c,
32'h5b865ba0,
32'h5bba5bd4,
32'h5bee5c08,
32'h5c225c3c,
32'h5c565c70,
32'h5c8a5ca4,
32'h5cbe5cd8,
32'h5cf25d0c,
32'h5d265d40,
32'h5d5a5d74,
32'h5d8e5da8,
32'h5dc25ddc,
32'h5df65e10,
32'h5e2a5e44,
32'h5e5e5e78,
32'h5e925eac,
32'h5ec65ee0,
32'h5efa5f14,
32'h5f2e5f48,
32'h5f625f7c,
32'h5f965fb0,
32'h5fca5fe4,
32'h5ffe6018,
32'h6032604c,
32'h60666080,
32'h60fe6118,
32'h6132614c,
32'h61666180,
32'h619a61b4,
32'h61ce61e8,
32'h6202621c,
32'h62366250,
32'h626a6284,
32'h629e62b8,
32'h62d262ec,
32'h63066320,
32'h633a6354,
32'h636e6388,
32'h63a263bc,
32'h63d663f0,
32'h640a6424,
32'h643e6458,
32'h6472648c,
32'h64a664c0,
32'h64da64f4,
32'h650e6528,
32'h6542655c,
32'h65766590,
32'h65aa65c4,
32'h65de65f8,
32'h6612662c,
32'h66466660,
32'h667a6694,
32'h66ae66c8,
32'h66e266fc,
32'h677a6794,
32'h67ae67c8,
32'h67e267fc,
32'h68166830,
32'h684a6864,
32'h687e6898,
32'h68b268cc,
32'h68e66900,
32'h691a6934,
32'h694e6968,
32'h6982699c,
32'h69b669d0,
32'h69ea6a04,
32'h6a1e6a38,
32'h6a526a6c,
32'h6a866aa0,
32'h6aba6ad4,
32'h6aee6b08,
32'h6b226b3c,
32'h6b566b70,
32'h6b8a6ba4,
32'h6bbe6bd8,
32'h6bf26c0c,
32'h6c266c40,
32'h6c5a6c74,
32'h6c8e6ca8,
32'h6cc26cdc,
32'h6cf66d10,
32'h6d2a6d44,
32'h6d5e6d78,
32'h6df66e10,
32'h6e2a6e44,
32'h6e5e6e78,
32'h6e926eac,
32'h6ec66ee0,
32'h6efa6f14,
32'h6f2e6f48,
32'h6f626f7c,
32'h6f966fb0,
32'h6fca6fe4,
32'h6ffe7018,
32'h7032704c,
32'h70667080,
32'h709a70b4,
32'h70ce70e8,
32'h7102711c,
32'h71367150,
32'h716a7184,
32'h719e71b8,
32'h71d271ec,
32'h72067220,
32'h723a7254,
32'h726e7288,
32'h72a272bc,
32'h72d672f0,
32'h730a7324,
32'h733e7358,
32'h7372738c,
32'h73a673c0,
32'h73da73f4,
32'h7472748c,
32'h74a674c0,
32'h74da74f4,
32'h750e7528,
32'h7542755c,
32'h75767590,
32'h75aa75c4,
32'h75de75f8,
32'h7612762c,
32'h76467660,
32'h767a7694,
32'h76ae76c8,
32'h76e276fc,
32'h77167730,
32'h774a7764,
32'h777e7798,
32'h77b277cc,
32'h77e67800,
32'h781a7834,
32'h784e7868,
32'h7882789c,
32'h78b678d0,
32'h78ea7904,
32'h791e7938,
32'h7952796c,
32'h798679a0,
32'h79ba79d4,
32'h79ee7a08,
32'h7a227a3c,
32'h7a567a70,
32'h7aee7b08,
32'h7b227b3c,
32'h7b567b70,
32'h7b8a7ba4,
32'h7bbe7bd8,
32'h7bf27c0c,
32'h7c267c40,
32'h7c5a7c74,
32'h7c8e7ca8,
32'h7cc27cdc,
32'h7cf67d10,
32'h7d2a7d44,
32'h7d5e7d78,
32'h7d927dac,
32'h7dc67de0,
32'h7dfa7e14,
32'h7e2e7e48,
32'h7e627e7c,
32'h7e967eb0,
32'h7eca7ee4,
32'h7efe7f18,
32'h7f327f4c,
32'h7f667f80,
32'h7f9a7fb4,
32'h7fce7fe8,
32'h8002801c,
32'h80368050,
32'h806a8084,
32'h809e80b8,
32'h80d280ec,
32'h816a8184,
32'h819e81b8,
32'h81d281ec,
32'h82068220,
32'h823a8254,
32'h826e8288,
32'h82a282bc,
32'h82d682f0,
32'h830a8324,
32'h833e8358,
32'h8372838c,
32'h83a683c0,
32'h83da83f4,
32'h840e8428,
32'h8442845c,
32'h84768490,
32'h84aa84c4,
32'h84de84f8,
32'h8512852c,
32'h85468560,
32'h857a8594,
32'h85ae85c8,
32'h85e285fc,
32'h86168630,
32'h864a8664,
32'h867e8698,
32'h86b286cc,
32'h86e68700,
32'h871a8734,
32'h874e8768,
32'h87e68800,
32'h881a8834,
32'h884e8868,
32'h8882889c,
32'h88b688d0,
32'h88ea8904,
32'h891e8938,
32'h8952896c,
32'h898689a0,
32'h89ba89d4,
32'h89ee8a08,
32'h8a228a3c,
32'h8a568a70,
32'h8a8a8aa4,
32'h8abe8ad8,
32'h8af28b0c,
32'h8b268b40,
32'h8b5a8b74,
32'h8b8e8ba8,
32'h8bc28bdc,
32'h8bf68c10,
32'h8c2a8c44,
32'h8c5e8c78,
32'h8c928cac,
32'h8cc68ce0,
32'h8cfa8d14,
32'h8d2e8d48,
32'h8d628d7c,
32'h8d968db0,
32'h8dca8de4,
32'h8e628e7c,
32'h8e968eb0,
32'h8eca8ee4,
32'h8efe8f18,
32'h8f328f4c,
32'h8f668f80,
32'h8f9a8fb4,
32'h8fce8fe8,
32'h9002901c,
32'h90369050,
32'h906a9084,
32'h909e90b8,
32'h90d290ec,
32'h91069120,
32'h913a9154,
32'h916e9188,
32'h91a291bc,
32'h91d691f0,
32'h920a9224,
32'h923e9258,
32'h9272928c,
32'h92a692c0,
32'h92da92f4,
32'h930e9328,
32'h9342935c,
32'h93769390,
32'h93aa93c4,
32'h93de93f8,
32'h9412942c,
32'h94469460,
32'h94de94f8,
32'h9512952c,
32'h95469560,
32'h957a9594,
32'h95ae95c8,
32'h95e295fc,
32'h96169630,
32'h964a9664,
32'h967e9698,
32'h96b296cc,
32'h96e69700,
32'h971a9734,
32'h974e9768,
32'h9782979c,
32'h97b697d0,
32'h97ea9804,
32'h981e9838,
32'h9852986c,
32'h988698a0,
32'h98ba98d4,
32'h98ee9908,
32'h9922993c,
32'h99569970,
32'h998a99a4,
32'h99be99d8,
32'h99f29a0c,
32'h9a269a40,
32'h9a5a9a74,
32'h9a8e9aa8,
32'h9ac29adc,
32'h9b5a9b74,
32'h9b8e9ba8,
32'h9bc29bdc,
32'h9bf69c10,
32'h9c2a9c44,
32'h9c5e9c78,
32'h9c929cac,
32'h9cc69ce0,
32'h9cfa9d14,
32'h9d2e9d48,
32'h9d629d7c,
32'h9d969db0,
32'h9dca9de4,
32'h9dfe9e18,
32'h9e329e4c,
32'h9e669e80,
32'h9e9a9eb4,
32'h9ece9ee8,
32'h9f029f1c,
32'h9f369f50,
32'h9f6a9f84,
32'h9f9e9fb8,
32'h9fd29fec,
32'ha006a020,
32'ha03aa054,
32'ha06ea088,
32'ha0a2a0bc,
32'ha0d6a0f0,
32'ha10aa124,
32'ha13ea158,
32'ha1d6a1f0,
32'ha20aa224,
32'ha23ea258,
32'ha272a28c,
32'ha2a6a2c0,
32'ha2daa2f4,
32'ha30ea328,
32'ha342a35c,
32'ha376a390,
32'ha3aaa3c4,
32'ha3dea3f8,
32'ha412a42c,
32'ha446a460,
32'ha47aa494,
32'ha4aea4c8,
32'ha4e2a4fc,
32'ha516a530,
32'ha54aa564,
32'ha57ea598,
32'ha5b2a5cc,
32'ha5e6a600,
32'ha61aa634,
32'ha64ea668,
32'ha682a69c,
32'ha6b6a6d0,
32'ha6eaa704,
32'ha71ea738,
32'ha752a76c,
32'ha786a7a0,
32'ha7baa7d4,
32'ha852a86c,
32'ha886a8a0,
32'ha8baa8d4,
32'ha8eea908,
32'ha922a93c,
32'ha956a970,
32'ha98aa9a4,
32'ha9bea9d8,
32'ha9f2aa0c,
32'haa26aa40,
32'haa5aaa74,
32'haa8eaaa8,
32'haac2aadc,
32'haaf6ab10,
32'hab2aab44,
32'hab5eab78,
32'hab92abac,
32'habc6abe0,
32'habfaac14,
32'hac2eac48,
32'hac62ac7c,
32'hac96acb0,
32'haccaace4,
32'hacfead18,
32'had32ad4c,
32'had66ad80,
32'had9aadb4,
32'hadceade8,
32'hae02ae1c,
32'hae36ae50,
32'haeceaee8,
32'haf02af1c,
32'haf36af50,
32'haf6aaf84,
32'haf9eafb8,
32'hafd2afec,
32'hb006b020,
32'hb03ab054,
32'hb06eb088,
32'hb0a2b0bc,
32'hb0d6b0f0,
32'hb10ab124,
32'hb13eb158,
32'hb172b18c,
32'hb1a6b1c0,
32'hb1dab1f4,
32'hb20eb228,
32'hb242b25c,
32'hb276b290,
32'hb2aab2c4,
32'hb2deb2f8,
32'hb312b32c,
32'hb346b360,
32'hb37ab394,
32'hb3aeb3c8,
32'hb3e2b3fc,
32'hb416b430,
32'hb44ab464,
32'hb47eb498,
32'hb4b2b4cc,
32'hb54ab564,
32'hb57eb598,
32'hb5b2b5cc,
32'hb5e6b600,
32'hb61ab634,
32'hb64eb668,
32'hb682b69c,
32'hb6b6b6d0,
32'hb6eab704,
32'hb71eb738,
32'hb752b76c,
32'hb786b7a0,
32'hb7bab7d4,
32'hb7eeb808,
32'hb822b83c,
32'hb856b870,
32'hb88ab8a4,
32'hb8beb8d8,
32'hb8f2b90c,
32'hb926b940,
32'hb95ab974,
32'hb98eb9a8,
32'hb9c2b9dc,
32'hb9f6ba10,
32'hba2aba44,
32'hba5eba78,
32'hba92baac,
32'hbac6bae0,
32'hbafabb14,
32'hbb2ebb48,
32'hbbc6bbe0,
32'hbbfabc14,
32'hbc2ebc48,
32'hbc62bc7c,
32'hbc96bcb0,
32'hbccabce4,
32'hbcfebd18,
32'hbd32bd4c,
32'hbd66bd80,
32'hbd9abdb4,
32'hbdcebde8,
32'hbe02be1c,
32'hbe36be50,
32'hbe6abe84,
32'hbe9ebeb8,
32'hbed2beec,
32'hbf06bf20,
32'hbf3abf54,
32'hbf6ebf88,
32'hbfa2bfbc,
32'hbfd6bff0,
32'hc00ac024,
32'hc03ec058,
32'hc072c08c,
32'hc0a6c0c0,
32'hc0dac0f4,
32'hc10ec128,
32'hc142c15c,
32'hc176c190,
32'hc1aac1c4
};
