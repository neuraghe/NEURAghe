// INSTRUCTION BUS PARAMETRES

// L2
`define NB_REGION 2

`define MASTER_0_REGION_0_START_ADDR 32'h1A00_0000
`define MASTER_0_REGION_0_END_ADDR   32'h1DFF_FFFF
`define MASTER_0_REGION_1_START_ADDR 32'h1C00_0000
`define MASTER_0_REGION_1_END_ADDR   32'h1FFF_FFFF
