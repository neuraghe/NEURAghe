VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO vbbgen_PULPV3_monitor
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN vbbgen_PULPV3_monitor 0 0 ;
  SIZE 85.85 BY 65.269 ;
  SYMMETRY X Y R90 ;
  PIN pwell_value_LB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.359 0 31.409 0.05 ;
    END
  END pwell_value_LB[0]
  PIN pwell_value_LB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.259 0 31.309 0.05 ;
    END
  END pwell_value_LB[1]
  PIN pwell_value_LB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.159 0 31.209 0.05 ;
    END
  END pwell_value_LB[2]
  PIN pwell_value_LB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.059 0 31.109 0.05 ;
    END
  END pwell_value_LB[3]
  PIN pwell_value_LB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.959 0 31.009 0.05 ;
    END
  END pwell_value_LB[4]
  PIN pwell_value_UB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.859 0 31.909 0.05 ;
    END
  END pwell_value_UB[0]
  PIN pwell_value_UB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.759 0 31.809 0.05 ;
    END
  END pwell_value_UB[1]
  PIN pwell_value_UB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.659 0 31.709 0.05 ;
    END
  END pwell_value_UB[2]
  PIN pwell_value_UB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.559 0 31.609 0.05 ;
    END
  END pwell_value_UB[3]
  PIN pwell_value_UB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 31.459 0 31.509 0.05 ;
    END
  END pwell_value_UB[4]
  PIN nwell_value_LB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.459 0 31.509 0.05 ;
    END
  END nwell_value_LB[0]
  PIN nwell_value_LB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.559 0 31.609 0.05 ;
    END
  END nwell_value_LB[1]
  PIN nwell_value_LB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.659 0 31.709 0.05 ;
    END
  END nwell_value_LB[2]
  PIN nwell_value_LB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.759 0 31.809 0.05 ;
    END
  END nwell_value_LB[3]
  PIN nwell_value_LB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.859 0 31.909 0.05 ;
    END
  END nwell_value_LB[4]
  PIN nwell_value_UB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.959 0 31.009 0.05 ;
    END
  END nwell_value_UB[0]
  PIN nwell_value_UB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.059 0 31.109 0.05 ;
    END
  END nwell_value_UB[1]
  PIN nwell_value_UB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.159 0 31.209 0.05 ;
    END
  END nwell_value_UB[2]
  PIN nwell_value_UB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.259 0 31.309 0.05 ;
    END
  END nwell_value_UB[3]
  PIN nwell_value_UB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.359 0 31.409 0.05 ;
    END
  END nwell_value_UB[4]
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 32.66 0.245 34.16 65.269 ;
        RECT 43.721 48.269 48.937 49.212 ;
        RECT 55.657 48.269 62.894 49.212 ;
        RECT 55.657 48.269 62.895 48.27 ;
        RECT 69.614 48.269 76.974 49.212 ;
        RECT 83.999 48.269 84.483 49.212 ;
      LAYER M4 ;
        RECT 85.613 3.165 85.723 63.508 ;
        RECT 0.691 63.007 85.723 63.117 ;
        RECT 85.389 3.165 85.723 63.117 ;
        RECT 31.741 62.783 85.723 63.117 ;
        RECT 58.915 3.333 85.723 3.533 ;
        RECT 57.649 0 59.55 0.11 ;
        RECT 58.915 0 59.249 3.6 ;
        RECT 42.872 65.159 44.142 65.269 ;
        RECT 43.233 62.783 43.567 65.269 ;
        RECT 0.691 48.621 32.13 49.021 ;
        RECT 18.98 8.209 30.651 8.459 ;
        RECT 18.98 12.28 30.627 12.53 ;
        RECT 0.724 23.866 30.081 24.2 ;
        RECT 18.98 18.068 29.759 18.318 ;
        RECT 18.98 22.132 29.338 22.382 ;
        RECT 0.724 25.45 29.103 25.784 ;
        RECT 18.98 7.716 19.23 24.2 ;
        RECT 13.76 7.716 19.23 7.966 ;
        RECT 13.76 6.526 14.203 6.636 ;
        RECT 14.093 6.411 14.203 6.636 ;
        RECT 13.76 6.526 14.01 7.966 ;
        RECT 0.691 43.086 13.05 43.42 ;
        RECT 1.331 48.486 1.523 49.021 ;
        RECT 0.691 65.159 1.259 65.269 ;
        RECT 0.691 43.086 1.091 62.893 ;
        RECT 0.724 23.866 1.058 62.893 ;
        RECT 0.691 43.086 0.801 65.269 ;
        RECT 83.999 48.269 84.483 49.212 ;
        RECT 69.756 48.269 76.974 49.212 ;
        RECT 43.863 48.269 48.795 49.212 ;
      LAYER M6 ;
        RECT 0 48.269 85.85 50.269 ;
      LAYER M3 ;
        RECT 44.87 48.609 75.919 48.859 ;
        RECT 75.669 48.142 75.919 48.859 ;
        RECT 44.87 33.166 45.12 48.859 ;
        RECT 31.826 33.166 45.12 33.416 ;
        RECT 29.792 8.209 32.13 8.459 ;
        RECT 30.15 12.28 32.13 12.53 ;
        RECT 27.988 12.292 28.205 12.5 ;
        RECT 27.988 18.106 28.205 18.314 ;
        RECT 27.698 12.292 27.916 12.5 ;
        RECT 27.698 18.106 27.916 18.314 ;
        RECT 20.916 12.292 21.134 12.5 ;
        RECT 20.916 18.106 21.134 18.314 ;
        RECT 20.627 12.292 20.844 12.5 ;
        RECT 20.627 18.106 20.844 18.314 ;
      LAYER M2 ;
        RECT 1.549 48.025 1.803 48.145 ;
        RECT 1.327 48.408 1.669 48.528 ;
        RECT 1.549 48.025 1.669 48.528 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.295 0 34.187 0.11 ;
    END
  END GND
  PIN VDD1V8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M3 ;
        RECT 18.98 7.314 19.23 15.431 ;
        RECT 13.674 7.314 19.23 7.498 ;
        RECT 13.674 2.5 13.858 7.498 ;
      LAYER M2 ;
        RECT 18.98 15.199 19.53 15.407 ;
        RECT 18.98 14.393 19.23 15.407 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.66 0.245 38.16 65.269 ;
        RECT 44.694 25.344 46.521 27.164 ;
      LAYER M4 ;
        RECT 44.711 25.344 46.504 27.164 ;
        RECT 33.883 3.82 37.779 4.12 ;
        RECT 33.883 9.227 37.779 9.527 ;
        RECT 33.883 14.689 37.779 14.989 ;
        RECT 33.883 20.116 37.779 20.416 ;
        RECT 33.883 25.561 37.779 25.861 ;
        RECT 33.883 30.031 37.779 30.331 ;
        RECT 33.883 38.621 37.779 38.921 ;
        RECT 33.883 44.055 37.779 44.355 ;
        RECT 33.883 50.09 37.779 50.39 ;
        RECT 33.883 56.688 37.779 56.988 ;
        RECT 33.883 62.13 37.779 62.43 ;
      LAYER M6 ;
        RECT 0 25.245 85.85 27.245 ;
      LAYER M3 ;
        RECT 29.405 31.513 46.605 32.513 ;
        RECT 44.605 17.019 46.605 32.513 ;
        RECT 29.405 26.616 30.405 32.513 ;
        RECT 18.525 28.272 30.405 28.522 ;
      LAYER M2 ;
        RECT 37.571 3.388 37.779 62.843 ;
        RECT 0 6.228 0.605 6.261 ;
        RECT 0 6.061 0.536 6.261 ;
        RECT 0.336 5.848 0.536 6.261 ;
        RECT 0 25.245 0.187 27.246 ;
        RECT 0 6.061 0.15 27.246 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.319 15.199 34.091 15.407 ;
    END
  END VDD1V8
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 29.242 20.961 30.807 21.169 ;
    END
    PORT
      LAYER M2 ;
        RECT 29.281 9.437 30.807 9.645 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.288 8.57 24.538 26.984 ;
        RECT 34.66 0.245 36.16 65.269 ;
      LAYER M6 ;
        RECT 0 10.245 85.85 12.245 ;
      LAYER M3 ;
        RECT 30.73 5.608 35.098 5.758 ;
        RECT 30.686 11.054 35.098 11.204 ;
        RECT 30.73 13.776 35.098 13.926 ;
        RECT 30.73 21.933 35.098 22.083 ;
        RECT 30.73 28.372 35.098 28.522 ;
        RECT 30.73 33.822 35.098 33.972 ;
        RECT 30.73 43.14 35.098 43.29 ;
        RECT 30.73 55.027 35.098 55.177 ;
        RECT 30.73 60.48 35.098 60.63 ;
        RECT 0.691 62.981 30.736 63.181 ;
        RECT 12.717 25.066 16.738 25.274 ;
        RECT 16.53 23.361 16.738 25.274 ;
        RECT 10.227 26.776 12.925 26.984 ;
        RECT 12.717 25.066 12.925 26.984 ;
        RECT 10.227 23.365 10.435 26.984 ;
        RECT 0.691 23.365 10.435 23.565 ;
        RECT 0.691 47.412 2.491 47.662 ;
        RECT 0.691 44.412 2.491 44.662 ;
        RECT 2.087 47.367 2.137 47.662 ;
        RECT 0.691 23.365 0.891 63.181 ;
        RECT 0.325 7.025 1.93 7.233 ;
        RECT 0.325 7.025 0.533 12.245 ;
      LAYER M2 ;
        RECT 0.691 23.361 30.807 23.569 ;
        RECT 29.416 10.648 30.707 11.873 ;
        RECT 12.047 25.066 21.337 25.274 ;
    END
    PORT
      LAYER M2 ;
        RECT 28.935 7.037 30.807 7.245 ;
    END
  END VDD
  PIN pwell_pos_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.291 0 0.341 0.05 ;
    END
  END pwell_pos_clk
  PIN pwell
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 5.182 2.761 13.867 3.211 ;
        RECT 13.417 2.761 13.867 7.493 ;
        RECT 13.417 7.043 23.174 7.493 ;
        RECT 22.724 7.043 23.174 28.179 ;
        RECT 22.724 27.729 29.013 28.179 ;
        RECT 28.563 27.729 29.013 46.891 ;
        RECT 28.563 46.441 30.388 46.891 ;
      LAYER M6 ;
        RECT 0 38.269 85.85 40.269 ;
    END
  END pwell
  PIN pwell_neg_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 32.059 0 32.109 0.05 ;
    END
  END pwell_neg_clk
  PIN compare_pwell_neg_LB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.859 0 30.909 0.05 ;
    END
  END compare_pwell_neg_LB
  PIN compare_pwell_neg_UB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 30.759 0 30.809 0.05 ;
    END
  END compare_pwell_neg_UB
  PIN compare_nwell_LB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.859 0 30.909 0.05 ;
    END
  END compare_nwell_LB
  PIN compare_nwell_UB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.759 0 30.809 0.05 ;
    END
  END compare_nwell_UB
  PIN nwell
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 29.871 13.225 30.239 17.245 ;
      LAYER M4 ;
        RECT 19.616 13.394 30.228 13.46 ;
      LAYER M6 ;
        RECT 0 15.245 85.85 17.245 ;
      LAYER M1 ;
        RECT 30.086 7.088 30.467 7.198 ;
        RECT 30.357 0.21 30.467 7.198 ;
        RECT 30.086 7.088 30.236 13.712 ;
    END
  END nwell
  PIN nwell_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 31.959 0 32.009 0.05 ;
    END
  END nwell_clk
  PIN compare_pwell_pos_LB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.659 0 30.709 0.05 ;
    END
  END compare_pwell_pos_LB
  PIN compare_pwell_pos_UB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 30.559 0 30.609 0.05 ;
    END
  END compare_pwell_pos_UB
  OBS
    LAYER M1 ;
      RECT 0 0 85.85 65.269 ;
    LAYER M2 ;
      RECT 0 0 85.85 65.269 ;
    LAYER M3 ;
      RECT 0 0 85.85 65.269 ;
    LAYER M4 ;
      RECT 0.033 25.278 0.167 27.212 ;
      RECT 0.291 0.55 0.341 6.933 ;
      RECT 0.362 10.278 0.496 12.212 ;
      RECT 1.697 43.873 1.847 44.049 ;
      RECT 1.747 43.853 1.797 46.722 ;
      RECT 1.432 25.937 9.806 32.711 ;
      RECT 1.432 32.923 11.406 42.897 ;
      RECT 3.075 6.526 13.26 6.776 ;
      RECT 0.696 0 13.87 1.974 ;
      RECT 1.353 49.647 14.527 62.821 ;
      RECT 10.031 26.649 15.986 26.983 ;
      RECT 14.503 24.303 14.623 24.671 ;
      RECT 14.503 24.605 17.8 24.671 ;
      RECT 0.696 8.42 13.26 23.194 ;
      RECT 0.696 8.466 18.48 23.194 ;
      RECT 15.116 24.371 20.752 24.437 ;
      RECT 21.605 17.844 21.861 17.894 ;
      RECT 19.516 17.146 22.463 17.212 ;
      RECT 24.288 22.493 24.538 23.569 ;
      RECT 24.288 20.491 24.538 22.021 ;
      RECT 24.288 18.453 24.538 20.205 ;
      RECT 24.288 10.401 24.538 12.153 ;
      RECT 24.288 8.57 24.538 10.114 ;
      RECT 12.301 26.213 12.415 26.413 ;
      RECT 12.301 26.363 25.966 26.413 ;
      RECT 27.365 22.55 27.415 22.806 ;
      RECT 27.365 7.8 27.415 8.056 ;
      RECT 14.745 49.647 27.919 62.821 ;
      RECT 19.352 20.315 29.316 20.381 ;
      RECT 19.352 20.315 19.462 20.736 ;
      RECT 19.354 12.979 29.316 13.045 ;
      RECT 19.354 12.979 19.42 14.629 ;
      RECT 19.516 10.225 29.316 10.291 ;
      RECT 19.516 10.225 19.668 10.738 ;
      RECT 1.353 47.921 30.384 48.321 ;
      RECT 29.603 25.45 30.386 25.784 ;
      RECT 9.969 24.941 30.386 25.275 ;
      RECT 14.093 0 30.467 5.911 ;
      RECT 14.703 0 30.467 6.774 ;
      RECT 30.559 0.55 30.609 6.931 ;
      RECT 18.644 6.881 30.609 6.931 ;
      RECT 30.659 0.55 30.709 7.081 ;
      RECT 18.64 7.031 30.709 7.081 ;
      RECT 30.284 24.31 30.763 24.376 ;
      RECT 30.284 24.31 30.35 24.837 ;
      RECT 19.516 17.561 30.763 17.627 ;
      RECT 30.759 0.55 30.809 7.231 ;
      RECT 30.859 0.55 30.909 7.381 ;
      RECT 30.959 0.55 31.009 24.275 ;
      RECT 31.059 0.55 31.109 23.22 ;
      RECT 31.159 0.55 31.209 23.823 ;
      RECT 31.259 0.55 31.309 20.593 ;
      RECT 31.359 0.55 31.409 18.414 ;
      RECT 31.459 0.55 31.509 15.137 ;
      RECT 31.559 0.55 31.609 12.974 ;
      RECT 31.659 0.55 31.709 10.254 ;
      RECT 31.759 0.55 31.809 7.293 ;
      RECT 31.859 0.55 31.909 23.53 ;
      RECT 31.959 0.55 32.009 24.516 ;
      RECT 30.473 24.466 32.009 24.516 ;
      RECT 30.473 24.466 30.587 24.658 ;
      RECT 32.059 0.55 32.109 46.992 ;
      RECT 39.281 61.611 39.615 62.345 ;
      RECT 38.6 49.253 38.75 62.611 ;
      RECT 40.682 62.007 40.832 62.611 ;
      RECT 38.6 62.461 40.832 62.611 ;
      RECT 1.301 63.617 42.733 64.659 ;
      RECT 1.759 63.617 42.372 65.269 ;
      RECT 34.687 0 57.149 2.934 ;
      RECT 32.282 0.61 58.415 2.934 ;
      RECT 63.139 62.007 63.289 62.611 ;
      RECT 63.139 3.619 63.289 4.222 ;
      RECT 63.439 4.045 63.589 4.648 ;
      RECT 84.881 50.62 85.215 50.754 ;
      RECT 85.065 50.62 85.215 53.312 ;
      RECT 85.065 12.917 85.215 15.609 ;
      RECT 84.881 15.475 85.215 15.609 ;
      RECT 44.067 63.617 85.113 64.659 ;
      RECT 44.642 64.008 85.723 65.269 ;
      RECT 60.05 0 85.85 2.665 ;
      RECT 59.749 0.61 84.889 2.833 ;
    LAYER M4 SPACING 0.05 ;
      RECT 0.033 25.278 0.167 27.212 ;
      RECT 0.362 10.278 0.496 12.212 ;
      RECT 0 62.985 0.584 65.269 ;
      RECT 0 63.288 0.599 65.269 ;
      RECT 0.998 23.672 10.12 23.774 ;
      RECT 0 0 0.199 23.774 ;
      RECT 0.433 0 13.87 1.974 ;
      RECT 0 0.142 13.668 2.393 ;
      RECT 0 6.526 13.668 6.776 ;
      RECT 0 0.142 13.567 6.918 ;
      RECT 0.291 0.142 0.341 6.933 ;
      RECT 0.64 7.34 13.567 23.258 ;
      RECT 0.64 7.605 13.668 23.258 ;
      RECT 0.64 8.279 18.888 8.389 ;
      RECT 0 0.142 0.218 23.774 ;
      RECT 0.64 8.058 18.873 23.254 ;
      RECT 2.037 0 13.567 23.258 ;
      RECT 0 12.352 16.423 23.258 ;
      RECT 0 12.352 0.584 23.774 ;
      RECT 10.542 8.058 16.423 23.774 ;
      RECT 16.845 15.538 18.888 23.774 ;
      RECT 29.438 26.663 30.372 27.197 ;
      RECT 34.712 60.488 35.046 60.622 ;
      RECT 34.712 55.035 35.046 55.169 ;
      RECT 34.712 43.148 35.046 43.282 ;
      RECT 34.712 33.83 35.046 33.964 ;
      RECT 34.712 28.38 35.046 28.514 ;
      RECT 34.712 21.941 35.046 22.075 ;
      RECT 34.712 13.784 35.046 13.918 ;
      RECT 34.712 11.062 35.046 11.196 ;
      RECT 34.712 5.616 35.046 5.75 ;
      RECT 37.013 31.633 37.807 32.393 ;
      RECT 30.843 63.209 43.141 65.067 ;
      RECT 0.893 63.288 43.141 65.067 ;
      RECT 1.351 63.288 42.78 65.269 ;
      RECT 14.093 0.142 32.203 5.501 ;
      RECT 63.139 3.619 63.289 62.691 ;
      RECT 14.093 0.202 58.823 3.728 ;
      RECT 34.279 0 57.557 3.728 ;
      RECT 14.093 0.202 33.791 5.501 ;
      RECT 14.093 4.212 85.297 5.501 ;
      RECT 14.093 0.142 30.709 6.319 ;
      RECT 30.759 0.142 30.809 8.102 ;
      RECT 30.859 0.142 30.909 8.102 ;
      RECT 31.759 0.142 31.809 8.102 ;
      RECT 14.093 0 30.467 6.319 ;
      RECT 14.295 0 30.467 7.207 ;
      RECT 14.102 6.728 85.297 7.207 ;
      RECT 19.337 5.865 85.297 8.102 ;
      RECT 19.337 0 29.685 8.117 ;
      RECT 31.659 0.142 31.709 10.947 ;
      RECT 32.237 5.865 85.297 9.135 ;
      RECT 35.205 4.212 85.297 9.135 ;
      RECT 19.337 8.566 33.791 10.947 ;
      RECT 19.337 9.619 85.297 10.947 ;
      RECT 19.337 8.566 30.579 12.173 ;
      RECT 19.337 11.311 85.297 12.173 ;
      RECT 19.337 8.551 29.685 12.185 ;
      RECT 19.337 8.551 20.52 12.188 ;
      RECT 21.241 8.551 27.591 12.188 ;
      RECT 28.312 8.566 30.043 12.188 ;
      RECT 19.337 12.622 30.043 13.302 ;
      RECT 31.559 0.142 31.609 13.669 ;
      RECT 19.337 12.637 85.297 13.302 ;
      RECT 19.337 12.622 19.524 17.976 ;
      RECT 30.32 12.637 85.297 13.669 ;
      RECT 32.237 11.311 85.297 13.669 ;
      RECT 19.337 13.552 30.623 15.092 ;
      RECT 35.205 9.619 85.297 14.597 ;
      RECT 19.337 14.033 85.297 14.597 ;
      RECT 19.337 14.033 33.791 15.092 ;
      RECT 31.459 0.142 31.509 15.137 ;
      RECT 19.337 13.552 28.212 17.976 ;
      RECT 31.259 0.142 31.309 21.826 ;
      RECT 31.359 0.142 31.409 21.826 ;
      RECT 31.496 14.033 31.546 21.826 ;
      RECT 37.871 0 57.557 16.912 ;
      RECT 19.337 15.514 44.498 17.976 ;
      RECT 19.322 15.538 44.498 17.976 ;
      RECT 19.322 18.41 20.52 22.04 ;
      RECT 21.241 18.41 27.591 22.04 ;
      RECT 29.851 15.514 44.498 20.024 ;
      RECT 34.198 15.081 44.498 20.024 ;
      RECT 19.322 18.421 33.791 21.826 ;
      RECT 19.322 20.508 44.498 21.826 ;
      RECT 28.312 18.41 30.763 22.04 ;
      RECT 19.322 18.421 30.763 22.04 ;
      RECT 30.959 0.142 31.009 28.265 ;
      RECT 31.059 0.142 31.109 28.265 ;
      RECT 31.159 0.142 31.209 28.265 ;
      RECT 31.859 0.142 31.909 28.265 ;
      RECT 31.959 0.142 32.009 28.265 ;
      RECT 29.43 18.41 30.763 23.774 ;
      RECT 19.322 22.474 44.498 23.774 ;
      RECT 30.173 22.19 44.498 25.469 ;
      RECT 10.542 24.371 44.498 24.437 ;
      RECT 10.542 24.605 44.498 24.671 ;
      RECT 10.542 24.292 16.423 25.275 ;
      RECT 1.15 24.941 44.498 25.275 ;
      RECT 1.15 24.292 10.12 25.358 ;
      RECT 10.542 24.292 12.61 25.358 ;
      RECT 16.845 24.292 44.498 25.358 ;
      RECT 35.205 20.508 44.498 25.469 ;
      RECT 29.195 24.292 33.791 26.509 ;
      RECT 10.542 26.363 44.498 26.413 ;
      RECT 10.542 25.876 12.61 26.983 ;
      RECT 1.15 26.649 29.298 26.983 ;
      RECT 1.15 25.876 10.12 42.994 ;
      RECT 13.032 25.876 29.298 28.165 ;
      RECT 1.15 27.854 44.498 27.92 ;
      RECT 30.512 25.953 44.498 28.265 ;
      RECT 1.15 28.234 30.386 28.568 ;
      RECT 30.512 15.514 30.623 31.406 ;
      RECT 35.205 25.953 44.498 29.939 ;
      RECT 30.512 28.629 44.498 29.939 ;
      RECT 30.512 28.629 33.791 31.406 ;
      RECT 37.871 0 44.498 31.406 ;
      RECT 30.512 30.423 44.498 31.406 ;
      RECT 1.15 28.629 29.298 42.994 ;
      RECT 46.712 3.692 85.297 48.035 ;
      RECT 1.15 32.62 85.297 33.059 ;
      RECT 1.15 32.62 31.719 33.715 ;
      RECT 1.15 33.523 44.763 33.715 ;
      RECT 1.15 27.091 18.418 42.994 ;
      RECT 35.205 33.523 44.763 38.529 ;
      RECT 1.15 34.079 44.763 38.529 ;
      RECT 1.15 34.079 33.791 42.994 ;
      RECT 13.142 39.013 44.763 43.033 ;
      RECT 13.142 32.62 30.623 48.529 ;
      RECT 32.059 0.142 32.109 48.529 ;
      RECT 13.142 43.397 44.763 43.963 ;
      RECT 35.205 39.013 44.763 43.963 ;
      RECT 1.183 43.512 33.791 44.305 ;
      RECT 1.747 43.512 1.797 47.305 ;
      RECT 1.183 44.769 44.763 47.26 ;
      RECT 1.183 44.769 1.98 47.305 ;
      RECT 2.244 44.769 44.763 47.305 ;
      RECT 2.598 43.512 33.791 48.529 ;
      RECT 59.341 3.625 85.297 48.035 ;
      RECT 37.871 33.523 44.763 48.177 ;
      RECT 45.227 32.62 75.562 48.177 ;
      RECT 76.026 3.625 85.297 48.177 ;
      RECT 1.183 47.769 43.771 48.394 ;
      RECT 48.887 3.692 69.664 48.502 ;
      RECT 1.183 47.769 1.239 48.529 ;
      RECT 1.615 47.769 43.771 48.529 ;
      RECT 49.147 0 49.447 62.691 ;
      RECT 49.747 0 50.047 62.691 ;
      RECT 50.347 0 50.647 62.691 ;
      RECT 50.947 0 51.247 62.691 ;
      RECT 51.547 0 51.847 62.691 ;
      RECT 52.147 0 52.447 62.691 ;
      RECT 52.747 0 53.047 62.691 ;
      RECT 53.347 0 53.647 62.691 ;
      RECT 53.947 0 54.247 62.691 ;
      RECT 54.547 0 54.847 62.691 ;
      RECT 55.147 0 55.447 62.691 ;
      RECT 55.799 3.692 62.753 62.691 ;
      RECT 63.104 3.625 63.404 62.691 ;
      RECT 63.704 3.625 64.004 62.691 ;
      RECT 64.304 3.625 64.604 62.691 ;
      RECT 64.904 3.625 65.204 62.691 ;
      RECT 65.504 3.625 65.804 62.691 ;
      RECT 66.104 3.625 66.404 62.691 ;
      RECT 66.704 3.625 67.004 62.691 ;
      RECT 67.304 3.625 67.604 62.691 ;
      RECT 67.904 3.625 68.204 62.691 ;
      RECT 68.504 3.625 68.804 62.691 ;
      RECT 69.104 3.625 69.404 62.691 ;
      RECT 48.887 48.966 69.664 62.691 ;
      RECT 77.066 3.625 83.907 62.691 ;
      RECT 32.222 44.447 43.771 49.998 ;
      RECT 1.183 49.113 33.791 54.92 ;
      RECT 1.183 50.482 85.297 54.92 ;
      RECT 35.205 50.482 85.297 56.596 ;
      RECT 1.183 55.284 85.297 56.596 ;
      RECT 1.183 55.284 33.791 60.373 ;
      RECT 1.183 57.08 85.297 60.373 ;
      RECT 1.183 49.113 30.623 62.874 ;
      RECT 35.205 57.08 85.297 62.038 ;
      RECT 1.183 60.737 85.297 62.038 ;
      RECT 1.183 60.737 33.791 62.691 ;
      RECT 37.871 49.304 85.297 62.691 ;
      RECT 84.575 3.625 85.297 62.691 ;
      RECT 1.183 62.522 85.297 62.691 ;
      RECT 1.183 60.737 31.649 62.874 ;
      RECT 30.843 60.737 31.649 62.915 ;
      RECT 43.659 63.209 85.521 65.067 ;
      RECT 44.234 63.6 85.85 65.269 ;
      RECT 59.642 0 85.85 3.073 ;
      RECT 59.341 0.202 85.297 3.241 ;
    LAYER M5 ;
      RECT 0.033 25.278 0.167 27.212 ;
      RECT 0.362 10.278 0.496 12.212 ;
      RECT 0.691 48.269 1.073 50.269 ;
      RECT 1.353 43.086 2.287 49.021 ;
      RECT 3.656 45.87 4.803 48.321 ;
      RECT 2.567 48.621 6.049 49.021 ;
      RECT 6.328 43.086 7.262 49.021 ;
      RECT 1.432 25.937 9.806 32.711 ;
      RECT 9.002 45.87 10.149 48.321 ;
      RECT 1.432 32.923 11.406 42.897 ;
      RECT 7.542 48.621 11.48 49.021 ;
      RECT 11.705 23.866 12.439 24.2 ;
      RECT 11.705 25.45 12.439 25.784 ;
      RECT 11.705 43.086 12.439 43.42 ;
      RECT 11.69 48.654 12.454 48.988 ;
      RECT 11.822 23.866 12.322 49.021 ;
      RECT 12.606 47.954 13.37 48.288 ;
      RECT 12.738 23.866 13.238 49.021 ;
      RECT 0.696 0 13.87 1.974 ;
      RECT 1.353 49.647 14.527 62.821 ;
      RECT 0.696 8.42 18.67 23.194 ;
      RECT 19.066 17.139 20.121 17.219 ;
      RECT 19.066 17.139 19.146 23.506 ;
      RECT 16.441 23.426 19.146 23.506 ;
      RECT 16.441 23.426 16.521 32.312 ;
      RECT 21.422 20.696 21.488 24.671 ;
      RECT 17.36 24.605 21.488 24.671 ;
      RECT 21.185 17.836 21.906 17.902 ;
      RECT 21.185 17.836 21.251 24.437 ;
      RECT 20.22 24.371 21.251 24.437 ;
      RECT 22.648 45.87 23.382 48.321 ;
      RECT 25.534 45.87 26.681 48.321 ;
      RECT 14.745 49.647 27.919 62.821 ;
      RECT 27.336 43.766 28.302 43.816 ;
      RECT 27.336 43.186 28.302 43.236 ;
      RECT 29.438 26.663 30.372 27.197 ;
      RECT 14.093 0 30.467 6.774 ;
      RECT 29.555 10.808 30.491 11.71 ;
      RECT 30.759 0.55 30.809 22.849 ;
      RECT 27.009 22.799 30.809 22.849 ;
      RECT 27.009 22.799 27.059 22.99 ;
      RECT 25.042 22.94 27.059 22.99 ;
      RECT 13.378 48.621 30.848 49.021 ;
      RECT 30.859 0.55 30.909 22.99 ;
      RECT 30.959 26.363 31.009 61.53 ;
      RECT 30.959 0.55 31.009 23.117 ;
      RECT 31.059 0.55 31.109 58.746 ;
      RECT 31.159 0.55 31.209 56.026 ;
      RECT 31.259 0.55 31.309 53.025 ;
      RECT 31.359 0.55 31.409 50.65 ;
      RECT 31.459 0.55 31.509 47.961 ;
      RECT 31.559 0.55 31.609 45.241 ;
      RECT 31.659 0.55 31.709 42.521 ;
      RECT 31.759 0.55 31.809 39.805 ;
      RECT 31.859 0.55 31.909 37.079 ;
      RECT 31.92 65.159 32.13 65.269 ;
      RECT 31.52 48.621 32.13 49.021 ;
      RECT 39.281 61.611 39.615 62.611 ;
      RECT 63.155 62.155 63.289 62.611 ;
      RECT 39.281 62.311 63.289 62.611 ;
      RECT 43.48 3.619 63.289 3.919 ;
      RECT 63.155 3.619 63.289 4.075 ;
      RECT 52.984 52.712 84.872 52.862 ;
      RECT 52.984 52.412 84.872 52.562 ;
      RECT 52.984 52.112 84.872 52.262 ;
      RECT 52.984 51.812 84.872 51.962 ;
      RECT 52.984 51.512 84.872 51.662 ;
      RECT 52.984 51.212 84.872 51.362 ;
      RECT 52.984 50.912 84.872 51.062 ;
      RECT 52.984 50.312 84.872 50.462 ;
      RECT 52.984 50.012 84.872 50.162 ;
      RECT 52.984 49.712 84.872 49.862 ;
      RECT 52.984 16.367 84.872 16.517 ;
      RECT 52.984 16.067 84.872 16.217 ;
      RECT 52.984 15.767 84.872 15.917 ;
      RECT 52.984 15.167 84.872 15.317 ;
      RECT 52.984 14.867 84.872 15.017 ;
      RECT 52.984 14.567 84.872 14.717 ;
      RECT 52.984 14.267 84.872 14.417 ;
      RECT 52.984 13.967 84.872 14.117 ;
      RECT 52.984 13.667 84.872 13.817 ;
      RECT 52.984 13.367 84.872 13.517 ;
      RECT 52.984 50.612 85.215 50.762 ;
      RECT 52.984 15.467 85.215 15.617 ;
    LAYER M5 SPACING 0.05 ;
      RECT 0.033 25.278 0.167 27.212 ;
      RECT 0 63 0.584 65.269 ;
      RECT 0.691 48.269 1.073 50.269 ;
      RECT 2.567 48.621 6.049 49.021 ;
      RECT 7.542 48.621 11.48 49.021 ;
      RECT 23.266 24.307 24.196 25.343 ;
      RECT 23.266 22.489 24.196 23.759 ;
      RECT 23.266 18.425 24.196 22.025 ;
      RECT 23.266 13.567 24.196 17.961 ;
      RECT 23.266 12.637 24.196 13.287 ;
      RECT 14.093 0 30.467 6.774 ;
      RECT 29.555 10.808 30.491 11.71 ;
      RECT 13.378 48.621 30.848 49.021 ;
      RECT 31.52 48.621 32.13 49.021 ;
      RECT 0.908 63.224 32.568 65.052 ;
      RECT 1.366 63.224 32.568 65.269 ;
      RECT 0 0 0.184 23.759 ;
      RECT 30.759 0.142 30.809 48.514 ;
      RECT 30.859 0.142 30.909 48.514 ;
      RECT 31.459 0.142 31.509 48.514 ;
      RECT 31.559 0.142 31.609 48.514 ;
      RECT 31.659 0.142 31.709 48.514 ;
      RECT 31.759 0.142 31.809 48.514 ;
      RECT 31.859 0.142 31.909 48.514 ;
      RECT 30.758 0.157 32.188 48.514 ;
      RECT 0.448 0 13.87 1.974 ;
      RECT 0 0.157 13.325 2.669 ;
      RECT 0 0.157 5.09 23.759 ;
      RECT 0 3.303 13.325 23.759 ;
      RECT 0 7.585 13.653 23.759 ;
      RECT 24.63 12.637 32.568 13.133 ;
      RECT 19.337 12.637 22.632 13.287 ;
      RECT 24.63 12.637 29.779 13.287 ;
      RECT 19.337 12.637 19.509 17.961 ;
      RECT 19.066 17.139 22.632 17.219 ;
      RECT 24.63 13.567 29.779 17.961 ;
      RECT 19.337 13.567 22.632 17.961 ;
      RECT 24.63 17.337 32.568 17.961 ;
      RECT 19.337 18.425 22.632 22.025 ;
      RECT 24.63 18.425 32.568 22.025 ;
      RECT 29.445 18.425 32.568 23.759 ;
      RECT 19.066 17.139 19.146 23.506 ;
      RECT 0 23.426 19.146 23.506 ;
      RECT 0 8.073 18.873 23.759 ;
      RECT 19.337 22.489 22.632 23.759 ;
      RECT 29.866 17.337 32.568 23.759 ;
      RECT 24.63 22.489 32.568 23.759 ;
      RECT 11.705 23.866 12.439 24.2 ;
      RECT 21.185 13.567 21.251 25.343 ;
      RECT 21.422 18.425 21.488 25.343 ;
      RECT 1.165 24.307 22.632 25.343 ;
      RECT 24.63 24.307 32.568 25.343 ;
      RECT 11.705 25.45 12.439 25.784 ;
      RECT 16.441 8.073 16.521 48.514 ;
      RECT 30.188 17.337 32.568 46.349 ;
      RECT 29.21 24.307 32.568 46.349 ;
      RECT 23.266 25.891 24.196 27.637 ;
      RECT 24.63 25.891 32.568 27.637 ;
      RECT 23.266 27.076 32.568 27.637 ;
      RECT 1.165 25.891 22.632 42.979 ;
      RECT 11.705 43.086 12.439 43.42 ;
      RECT 12.738 28.271 28.471 48.514 ;
      RECT 30.331 12.637 32.568 46.349 ;
      RECT 29.105 25.891 32.568 46.349 ;
      RECT 30.734 8.566 32.568 48.514 ;
      RECT 30.48 12.637 32.568 48.514 ;
      RECT 1.198 43.527 28.471 48.379 ;
      RECT 30.758 0.217 32.568 48.514 ;
      RECT 1.353 46.983 32.568 48.514 ;
      RECT 11.69 48.654 12.454 48.988 ;
      RECT 1.353 43.086 2.287 49.021 ;
      RECT 6.328 43.086 7.262 49.021 ;
      RECT 11.822 23.866 12.322 49.021 ;
      RECT 12.738 23.866 13.238 49.021 ;
      RECT 30.959 0.142 31.009 62.9 ;
      RECT 31.059 0.142 31.109 62.9 ;
      RECT 31.159 0.142 31.209 62.9 ;
      RECT 31.259 0.142 31.309 62.9 ;
      RECT 31.359 0.142 31.409 62.9 ;
      RECT 32.237 0.217 32.568 62.676 ;
      RECT 1.198 49.128 32.568 62.676 ;
      RECT 1.198 49.128 31.634 62.9 ;
      RECT 34.252 30.438 34.568 38.514 ;
      RECT 36.252 30.438 36.568 38.514 ;
      RECT 38.252 63.224 43.126 65.052 ;
      RECT 38.252 63.224 42.765 65.269 ;
      RECT 37.886 0 57.542 0.153 ;
      RECT 38.252 0.217 58.808 25.237 ;
      RECT 38.252 3.619 63.289 25.237 ;
      RECT 38.252 0 57.542 25.237 ;
      RECT 38.252 0 44.604 25.252 ;
      RECT 46.611 3.64 85.282 25.252 ;
      RECT 38.252 0 44.602 48.162 ;
      RECT 38.252 27.256 44.604 48.162 ;
      RECT 46.611 27.256 85.282 48.162 ;
      RECT 46.613 3.64 85.282 48.162 ;
      RECT 38.252 27.271 85.282 48.162 ;
      RECT 38.252 0 43.756 48.177 ;
      RECT 48.902 3.64 69.649 48.177 ;
      RECT 38.252 0 43.629 62.676 ;
      RECT 49.029 0 55.565 62.676 ;
      RECT 62.987 3.64 69.522 62.676 ;
      RECT 62.986 48.362 69.522 62.676 ;
      RECT 38.252 49.304 43.756 62.676 ;
      RECT 48.902 49.304 69.649 62.676 ;
      RECT 77.066 48.269 77.23 62.676 ;
      RECT 76.974 49.304 77.23 62.676 ;
      RECT 38.252 49.319 85.282 62.676 ;
      RECT 43.674 63.224 85.506 65.052 ;
      RECT 44.249 63.615 85.85 65.269 ;
      RECT 59.657 0 85.85 3.058 ;
      RECT 59.356 0.217 85.282 3.226 ;
  END
END vbbgen_PULPV3_monitor

END LIBRARY
