task ddr_x_readmem_32x8_ramloops;
  $readmemh("slm_files/ddr_x_mem_cut0_0.slm", `DDR_X_BRAM_RAMLOOP(0) );
  $readmemh("slm_files/ddr_x_mem_cut1_0.slm", `DDR_X_BRAM_RAMLOOP(1) );
  $readmemh("slm_files/ddr_x_mem_cut2_0.slm", `DDR_X_BRAM_RAMLOOP(2) );
  $readmemh("slm_files/ddr_x_mem_cut3_0.slm", `DDR_X_BRAM_RAMLOOP(3) );
  $readmemh("slm_files/ddr_x_mem_cut4_0.slm", `DDR_X_BRAM_RAMLOOP(4) );
  $readmemh("slm_files/ddr_x_mem_cut5_0.slm", `DDR_X_BRAM_RAMLOOP(5) );
  $readmemh("slm_files/ddr_x_mem_cut6_0.slm", `DDR_X_BRAM_RAMLOOP(6) );
  $readmemh("slm_files/ddr_x_mem_cut7_0.slm", `DDR_X_BRAM_RAMLOOP(7) );
  $readmemh("slm_files/ddr_x_mem_cut8_0.slm", `DDR_X_BRAM_RAMLOOP(8) );
  $readmemh("slm_files/ddr_x_mem_cut9_0.slm", `DDR_X_BRAM_RAMLOOP(9) );
  $readmemh("slm_files/ddr_x_mem_cut10_0.slm", `DDR_X_BRAM_RAMLOOP(10) );
  $readmemh("slm_files/ddr_x_mem_cut11_0.slm", `DDR_X_BRAM_RAMLOOP(11) );
  $readmemh("slm_files/ddr_x_mem_cut12_0.slm", `DDR_X_BRAM_RAMLOOP(12) );
  $readmemh("slm_files/ddr_x_mem_cut13_0.slm", `DDR_X_BRAM_RAMLOOP(13) );
  $readmemh("slm_files/ddr_x_mem_cut14_0.slm", `DDR_X_BRAM_RAMLOOP(14) );
  $readmemh("slm_files/ddr_x_mem_cut15_0.slm", `DDR_X_BRAM_RAMLOOP(15) );
  $readmemh("slm_files/ddr_x_mem_cut16_0.slm", `DDR_X_BRAM_RAMLOOP(16) );
  $readmemh("slm_files/ddr_x_mem_cut17_0.slm", `DDR_X_BRAM_RAMLOOP(17) );
  $readmemh("slm_files/ddr_x_mem_cut18_0.slm", `DDR_X_BRAM_RAMLOOP(18) );
  $readmemh("slm_files/ddr_x_mem_cut19_0.slm", `DDR_X_BRAM_RAMLOOP(19) );
  $readmemh("slm_files/ddr_x_mem_cut20_0.slm", `DDR_X_BRAM_RAMLOOP(20) );
  $readmemh("slm_files/ddr_x_mem_cut21_0.slm", `DDR_X_BRAM_RAMLOOP(21) );
  $readmemh("slm_files/ddr_x_mem_cut22_0.slm", `DDR_X_BRAM_RAMLOOP(22) );
  $readmemh("slm_files/ddr_x_mem_cut23_0.slm", `DDR_X_BRAM_RAMLOOP(23) );
  $readmemh("slm_files/ddr_x_mem_cut24_0.slm", `DDR_X_BRAM_RAMLOOP(24) );
  $readmemh("slm_files/ddr_x_mem_cut25_0.slm", `DDR_X_BRAM_RAMLOOP(25) );
  $readmemh("slm_files/ddr_x_mem_cut26_0.slm", `DDR_X_BRAM_RAMLOOP(26) );
  $readmemh("slm_files/ddr_x_mem_cut27_0.slm", `DDR_X_BRAM_RAMLOOP(27) );
  $readmemh("slm_files/ddr_x_mem_cut28_0.slm", `DDR_X_BRAM_RAMLOOP(28) );
  $readmemh("slm_files/ddr_x_mem_cut29_0.slm", `DDR_X_BRAM_RAMLOOP(29) );
  $readmemh("slm_files/ddr_x_mem_cut30_0.slm", `DDR_X_BRAM_RAMLOOP(30) );
  $readmemh("slm_files/ddr_x_mem_cut31_0.slm", `DDR_X_BRAM_RAMLOOP(31) );
  $readmemh("slm_files/ddr_x_mem_cut0_1.slm", `DDR_X_BRAM_RAMLOOP(32) );
  $readmemh("slm_files/ddr_x_mem_cut1_1.slm", `DDR_X_BRAM_RAMLOOP(33) );
  $readmemh("slm_files/ddr_x_mem_cut2_1.slm", `DDR_X_BRAM_RAMLOOP(34) );
  $readmemh("slm_files/ddr_x_mem_cut3_1.slm", `DDR_X_BRAM_RAMLOOP(35) );
  $readmemh("slm_files/ddr_x_mem_cut4_1.slm", `DDR_X_BRAM_RAMLOOP(36) );
  $readmemh("slm_files/ddr_x_mem_cut5_1.slm", `DDR_X_BRAM_RAMLOOP(37) );
  $readmemh("slm_files/ddr_x_mem_cut6_1.slm", `DDR_X_BRAM_RAMLOOP(38) );
  $readmemh("slm_files/ddr_x_mem_cut7_1.slm", `DDR_X_BRAM_RAMLOOP(39) );
  $readmemh("slm_files/ddr_x_mem_cut8_1.slm", `DDR_X_BRAM_RAMLOOP(40) );
  $readmemh("slm_files/ddr_x_mem_cut9_1.slm", `DDR_X_BRAM_RAMLOOP(41) );
  $readmemh("slm_files/ddr_x_mem_cut10_1.slm", `DDR_X_BRAM_RAMLOOP(42) );
  $readmemh("slm_files/ddr_x_mem_cut11_1.slm", `DDR_X_BRAM_RAMLOOP(43) );
  $readmemh("slm_files/ddr_x_mem_cut12_1.slm", `DDR_X_BRAM_RAMLOOP(44) );
  $readmemh("slm_files/ddr_x_mem_cut13_1.slm", `DDR_X_BRAM_RAMLOOP(45) );
  $readmemh("slm_files/ddr_x_mem_cut14_1.slm", `DDR_X_BRAM_RAMLOOP(46) );
  $readmemh("slm_files/ddr_x_mem_cut15_1.slm", `DDR_X_BRAM_RAMLOOP(47) );
  $readmemh("slm_files/ddr_x_mem_cut16_1.slm", `DDR_X_BRAM_RAMLOOP(48) );
  $readmemh("slm_files/ddr_x_mem_cut17_1.slm", `DDR_X_BRAM_RAMLOOP(49) );
  $readmemh("slm_files/ddr_x_mem_cut18_1.slm", `DDR_X_BRAM_RAMLOOP(50) );
  $readmemh("slm_files/ddr_x_mem_cut19_1.slm", `DDR_X_BRAM_RAMLOOP(51) );
  $readmemh("slm_files/ddr_x_mem_cut20_1.slm", `DDR_X_BRAM_RAMLOOP(52) );
  $readmemh("slm_files/ddr_x_mem_cut21_1.slm", `DDR_X_BRAM_RAMLOOP(53) );
  $readmemh("slm_files/ddr_x_mem_cut22_1.slm", `DDR_X_BRAM_RAMLOOP(54) );
  $readmemh("slm_files/ddr_x_mem_cut23_1.slm", `DDR_X_BRAM_RAMLOOP(55) );
  $readmemh("slm_files/ddr_x_mem_cut24_1.slm", `DDR_X_BRAM_RAMLOOP(56) );
  $readmemh("slm_files/ddr_x_mem_cut25_1.slm", `DDR_X_BRAM_RAMLOOP(57) );
  $readmemh("slm_files/ddr_x_mem_cut26_1.slm", `DDR_X_BRAM_RAMLOOP(58) );
  $readmemh("slm_files/ddr_x_mem_cut27_1.slm", `DDR_X_BRAM_RAMLOOP(59) );
  $readmemh("slm_files/ddr_x_mem_cut28_1.slm", `DDR_X_BRAM_RAMLOOP(60) );
  $readmemh("slm_files/ddr_x_mem_cut29_1.slm", `DDR_X_BRAM_RAMLOOP(61) );
  $readmemh("slm_files/ddr_x_mem_cut30_1.slm", `DDR_X_BRAM_RAMLOOP(62) );
  $readmemh("slm_files/ddr_x_mem_cut31_1.slm", `DDR_X_BRAM_RAMLOOP(63) );
  $readmemh("slm_files/ddr_x_mem_cut0_2.slm", `DDR_X_BRAM_RAMLOOP(64) );
  $readmemh("slm_files/ddr_x_mem_cut1_2.slm", `DDR_X_BRAM_RAMLOOP(65) );
  $readmemh("slm_files/ddr_x_mem_cut2_2.slm", `DDR_X_BRAM_RAMLOOP(66) );
  $readmemh("slm_files/ddr_x_mem_cut3_2.slm", `DDR_X_BRAM_RAMLOOP(67) );
  $readmemh("slm_files/ddr_x_mem_cut4_2.slm", `DDR_X_BRAM_RAMLOOP(68) );
  $readmemh("slm_files/ddr_x_mem_cut5_2.slm", `DDR_X_BRAM_RAMLOOP(69) );
  $readmemh("slm_files/ddr_x_mem_cut6_2.slm", `DDR_X_BRAM_RAMLOOP(70) );
  $readmemh("slm_files/ddr_x_mem_cut7_2.slm", `DDR_X_BRAM_RAMLOOP(71) );
  $readmemh("slm_files/ddr_x_mem_cut8_2.slm", `DDR_X_BRAM_RAMLOOP(72) );
  $readmemh("slm_files/ddr_x_mem_cut9_2.slm", `DDR_X_BRAM_RAMLOOP(73) );
  $readmemh("slm_files/ddr_x_mem_cut10_2.slm", `DDR_X_BRAM_RAMLOOP(74) );
  $readmemh("slm_files/ddr_x_mem_cut11_2.slm", `DDR_X_BRAM_RAMLOOP(75) );
  $readmemh("slm_files/ddr_x_mem_cut12_2.slm", `DDR_X_BRAM_RAMLOOP(76) );
  $readmemh("slm_files/ddr_x_mem_cut13_2.slm", `DDR_X_BRAM_RAMLOOP(77) );
  $readmemh("slm_files/ddr_x_mem_cut14_2.slm", `DDR_X_BRAM_RAMLOOP(78) );
  $readmemh("slm_files/ddr_x_mem_cut15_2.slm", `DDR_X_BRAM_RAMLOOP(79) );
  $readmemh("slm_files/ddr_x_mem_cut16_2.slm", `DDR_X_BRAM_RAMLOOP(80) );
  $readmemh("slm_files/ddr_x_mem_cut17_2.slm", `DDR_X_BRAM_RAMLOOP(81) );
  $readmemh("slm_files/ddr_x_mem_cut18_2.slm", `DDR_X_BRAM_RAMLOOP(82) );
  $readmemh("slm_files/ddr_x_mem_cut19_2.slm", `DDR_X_BRAM_RAMLOOP(83) );
  $readmemh("slm_files/ddr_x_mem_cut20_2.slm", `DDR_X_BRAM_RAMLOOP(84) );
  $readmemh("slm_files/ddr_x_mem_cut21_2.slm", `DDR_X_BRAM_RAMLOOP(85) );
  $readmemh("slm_files/ddr_x_mem_cut22_2.slm", `DDR_X_BRAM_RAMLOOP(86) );
  $readmemh("slm_files/ddr_x_mem_cut23_2.slm", `DDR_X_BRAM_RAMLOOP(87) );
  $readmemh("slm_files/ddr_x_mem_cut24_2.slm", `DDR_X_BRAM_RAMLOOP(88) );
  $readmemh("slm_files/ddr_x_mem_cut25_2.slm", `DDR_X_BRAM_RAMLOOP(89) );
  $readmemh("slm_files/ddr_x_mem_cut26_2.slm", `DDR_X_BRAM_RAMLOOP(90) );
  $readmemh("slm_files/ddr_x_mem_cut27_2.slm", `DDR_X_BRAM_RAMLOOP(91) );
  $readmemh("slm_files/ddr_x_mem_cut28_2.slm", `DDR_X_BRAM_RAMLOOP(92) );
  $readmemh("slm_files/ddr_x_mem_cut29_2.slm", `DDR_X_BRAM_RAMLOOP(93) );
  $readmemh("slm_files/ddr_x_mem_cut30_2.slm", `DDR_X_BRAM_RAMLOOP(94) );
  $readmemh("slm_files/ddr_x_mem_cut31_2.slm", `DDR_X_BRAM_RAMLOOP(95) );
  $readmemh("slm_files/ddr_x_mem_cut0_3.slm", `DDR_X_BRAM_RAMLOOP(96) );
  $readmemh("slm_files/ddr_x_mem_cut1_3.slm", `DDR_X_BRAM_RAMLOOP(97) );
  $readmemh("slm_files/ddr_x_mem_cut2_3.slm", `DDR_X_BRAM_RAMLOOP(98) );
  $readmemh("slm_files/ddr_x_mem_cut3_3.slm", `DDR_X_BRAM_RAMLOOP(99) );
  $readmemh("slm_files/ddr_x_mem_cut4_3.slm", `DDR_X_BRAM_RAMLOOP(100) );
  $readmemh("slm_files/ddr_x_mem_cut5_3.slm", `DDR_X_BRAM_RAMLOOP(101) );
  $readmemh("slm_files/ddr_x_mem_cut6_3.slm", `DDR_X_BRAM_RAMLOOP(102) );
  $readmemh("slm_files/ddr_x_mem_cut7_3.slm", `DDR_X_BRAM_RAMLOOP(103) );
  $readmemh("slm_files/ddr_x_mem_cut8_3.slm", `DDR_X_BRAM_RAMLOOP(104) );
  $readmemh("slm_files/ddr_x_mem_cut9_3.slm", `DDR_X_BRAM_RAMLOOP(105) );
  $readmemh("slm_files/ddr_x_mem_cut10_3.slm", `DDR_X_BRAM_RAMLOOP(106) );
  $readmemh("slm_files/ddr_x_mem_cut11_3.slm", `DDR_X_BRAM_RAMLOOP(107) );
  $readmemh("slm_files/ddr_x_mem_cut12_3.slm", `DDR_X_BRAM_RAMLOOP(108) );
  $readmemh("slm_files/ddr_x_mem_cut13_3.slm", `DDR_X_BRAM_RAMLOOP(109) );
  $readmemh("slm_files/ddr_x_mem_cut14_3.slm", `DDR_X_BRAM_RAMLOOP(110) );
  $readmemh("slm_files/ddr_x_mem_cut15_3.slm", `DDR_X_BRAM_RAMLOOP(111) );
  $readmemh("slm_files/ddr_x_mem_cut16_3.slm", `DDR_X_BRAM_RAMLOOP(112) );
  $readmemh("slm_files/ddr_x_mem_cut17_3.slm", `DDR_X_BRAM_RAMLOOP(113) );
  $readmemh("slm_files/ddr_x_mem_cut18_3.slm", `DDR_X_BRAM_RAMLOOP(114) );
  $readmemh("slm_files/ddr_x_mem_cut19_3.slm", `DDR_X_BRAM_RAMLOOP(115) );
  $readmemh("slm_files/ddr_x_mem_cut20_3.slm", `DDR_X_BRAM_RAMLOOP(116) );
  $readmemh("slm_files/ddr_x_mem_cut21_3.slm", `DDR_X_BRAM_RAMLOOP(117) );
  $readmemh("slm_files/ddr_x_mem_cut22_3.slm", `DDR_X_BRAM_RAMLOOP(118) );
  $readmemh("slm_files/ddr_x_mem_cut23_3.slm", `DDR_X_BRAM_RAMLOOP(119) );
  $readmemh("slm_files/ddr_x_mem_cut24_3.slm", `DDR_X_BRAM_RAMLOOP(120) );
  $readmemh("slm_files/ddr_x_mem_cut25_3.slm", `DDR_X_BRAM_RAMLOOP(121) );
  $readmemh("slm_files/ddr_x_mem_cut26_3.slm", `DDR_X_BRAM_RAMLOOP(122) );
  $readmemh("slm_files/ddr_x_mem_cut27_3.slm", `DDR_X_BRAM_RAMLOOP(123) );
  $readmemh("slm_files/ddr_x_mem_cut28_3.slm", `DDR_X_BRAM_RAMLOOP(124) );
  $readmemh("slm_files/ddr_x_mem_cut29_3.slm", `DDR_X_BRAM_RAMLOOP(125) );
  $readmemh("slm_files/ddr_x_mem_cut30_3.slm", `DDR_X_BRAM_RAMLOOP(126) );
  $readmemh("slm_files/ddr_x_mem_cut31_3.slm", `DDR_X_BRAM_RAMLOOP(127) );
  $readmemh("slm_files/ddr_x_mem_cut0_4.slm", `DDR_X_BRAM_RAMLOOP(128) );
  $readmemh("slm_files/ddr_x_mem_cut1_4.slm", `DDR_X_BRAM_RAMLOOP(129) );
  $readmemh("slm_files/ddr_x_mem_cut2_4.slm", `DDR_X_BRAM_RAMLOOP(130) );
  $readmemh("slm_files/ddr_x_mem_cut3_4.slm", `DDR_X_BRAM_RAMLOOP(131) );
  $readmemh("slm_files/ddr_x_mem_cut4_4.slm", `DDR_X_BRAM_RAMLOOP(132) );
  $readmemh("slm_files/ddr_x_mem_cut5_4.slm", `DDR_X_BRAM_RAMLOOP(133) );
  $readmemh("slm_files/ddr_x_mem_cut6_4.slm", `DDR_X_BRAM_RAMLOOP(134) );
  $readmemh("slm_files/ddr_x_mem_cut7_4.slm", `DDR_X_BRAM_RAMLOOP(135) );
  $readmemh("slm_files/ddr_x_mem_cut8_4.slm", `DDR_X_BRAM_RAMLOOP(136) );
  $readmemh("slm_files/ddr_x_mem_cut9_4.slm", `DDR_X_BRAM_RAMLOOP(137) );
  $readmemh("slm_files/ddr_x_mem_cut10_4.slm", `DDR_X_BRAM_RAMLOOP(138) );
  $readmemh("slm_files/ddr_x_mem_cut11_4.slm", `DDR_X_BRAM_RAMLOOP(139) );
  $readmemh("slm_files/ddr_x_mem_cut12_4.slm", `DDR_X_BRAM_RAMLOOP(140) );
  $readmemh("slm_files/ddr_x_mem_cut13_4.slm", `DDR_X_BRAM_RAMLOOP(141) );
  $readmemh("slm_files/ddr_x_mem_cut14_4.slm", `DDR_X_BRAM_RAMLOOP(142) );
  $readmemh("slm_files/ddr_x_mem_cut15_4.slm", `DDR_X_BRAM_RAMLOOP(143) );
  $readmemh("slm_files/ddr_x_mem_cut16_4.slm", `DDR_X_BRAM_RAMLOOP(144) );
  $readmemh("slm_files/ddr_x_mem_cut17_4.slm", `DDR_X_BRAM_RAMLOOP(145) );
  $readmemh("slm_files/ddr_x_mem_cut18_4.slm", `DDR_X_BRAM_RAMLOOP(146) );
  $readmemh("slm_files/ddr_x_mem_cut19_4.slm", `DDR_X_BRAM_RAMLOOP(147) );
  $readmemh("slm_files/ddr_x_mem_cut20_4.slm", `DDR_X_BRAM_RAMLOOP(148) );
  $readmemh("slm_files/ddr_x_mem_cut21_4.slm", `DDR_X_BRAM_RAMLOOP(149) );
  $readmemh("slm_files/ddr_x_mem_cut22_4.slm", `DDR_X_BRAM_RAMLOOP(150) );
  $readmemh("slm_files/ddr_x_mem_cut23_4.slm", `DDR_X_BRAM_RAMLOOP(151) );
  $readmemh("slm_files/ddr_x_mem_cut24_4.slm", `DDR_X_BRAM_RAMLOOP(152) );
  $readmemh("slm_files/ddr_x_mem_cut25_4.slm", `DDR_X_BRAM_RAMLOOP(153) );
  $readmemh("slm_files/ddr_x_mem_cut26_4.slm", `DDR_X_BRAM_RAMLOOP(154) );
  $readmemh("slm_files/ddr_x_mem_cut27_4.slm", `DDR_X_BRAM_RAMLOOP(155) );
  $readmemh("slm_files/ddr_x_mem_cut28_4.slm", `DDR_X_BRAM_RAMLOOP(156) );
  $readmemh("slm_files/ddr_x_mem_cut29_4.slm", `DDR_X_BRAM_RAMLOOP(157) );
  $readmemh("slm_files/ddr_x_mem_cut30_4.slm", `DDR_X_BRAM_RAMLOOP(158) );
  $readmemh("slm_files/ddr_x_mem_cut31_4.slm", `DDR_X_BRAM_RAMLOOP(159) );
  $readmemh("slm_files/ddr_x_mem_cut0_5.slm", `DDR_X_BRAM_RAMLOOP(160) );
  $readmemh("slm_files/ddr_x_mem_cut1_5.slm", `DDR_X_BRAM_RAMLOOP(161) );
  $readmemh("slm_files/ddr_x_mem_cut2_5.slm", `DDR_X_BRAM_RAMLOOP(162) );
  $readmemh("slm_files/ddr_x_mem_cut3_5.slm", `DDR_X_BRAM_RAMLOOP(163) );
  $readmemh("slm_files/ddr_x_mem_cut4_5.slm", `DDR_X_BRAM_RAMLOOP(164) );
  $readmemh("slm_files/ddr_x_mem_cut5_5.slm", `DDR_X_BRAM_RAMLOOP(165) );
  $readmemh("slm_files/ddr_x_mem_cut6_5.slm", `DDR_X_BRAM_RAMLOOP(166) );
  $readmemh("slm_files/ddr_x_mem_cut7_5.slm", `DDR_X_BRAM_RAMLOOP(167) );
  $readmemh("slm_files/ddr_x_mem_cut8_5.slm", `DDR_X_BRAM_RAMLOOP(168) );
  $readmemh("slm_files/ddr_x_mem_cut9_5.slm", `DDR_X_BRAM_RAMLOOP(169) );
  $readmemh("slm_files/ddr_x_mem_cut10_5.slm", `DDR_X_BRAM_RAMLOOP(170) );
  $readmemh("slm_files/ddr_x_mem_cut11_5.slm", `DDR_X_BRAM_RAMLOOP(171) );
  $readmemh("slm_files/ddr_x_mem_cut12_5.slm", `DDR_X_BRAM_RAMLOOP(172) );
  $readmemh("slm_files/ddr_x_mem_cut13_5.slm", `DDR_X_BRAM_RAMLOOP(173) );
  $readmemh("slm_files/ddr_x_mem_cut14_5.slm", `DDR_X_BRAM_RAMLOOP(174) );
  $readmemh("slm_files/ddr_x_mem_cut15_5.slm", `DDR_X_BRAM_RAMLOOP(175) );
  $readmemh("slm_files/ddr_x_mem_cut16_5.slm", `DDR_X_BRAM_RAMLOOP(176) );
  $readmemh("slm_files/ddr_x_mem_cut17_5.slm", `DDR_X_BRAM_RAMLOOP(177) );
  $readmemh("slm_files/ddr_x_mem_cut18_5.slm", `DDR_X_BRAM_RAMLOOP(178) );
  $readmemh("slm_files/ddr_x_mem_cut19_5.slm", `DDR_X_BRAM_RAMLOOP(179) );
  $readmemh("slm_files/ddr_x_mem_cut20_5.slm", `DDR_X_BRAM_RAMLOOP(180) );
  $readmemh("slm_files/ddr_x_mem_cut21_5.slm", `DDR_X_BRAM_RAMLOOP(181) );
  $readmemh("slm_files/ddr_x_mem_cut22_5.slm", `DDR_X_BRAM_RAMLOOP(182) );
  $readmemh("slm_files/ddr_x_mem_cut23_5.slm", `DDR_X_BRAM_RAMLOOP(183) );
  $readmemh("slm_files/ddr_x_mem_cut24_5.slm", `DDR_X_BRAM_RAMLOOP(184) );
  $readmemh("slm_files/ddr_x_mem_cut25_5.slm", `DDR_X_BRAM_RAMLOOP(185) );
  $readmemh("slm_files/ddr_x_mem_cut26_5.slm", `DDR_X_BRAM_RAMLOOP(186) );
  $readmemh("slm_files/ddr_x_mem_cut27_5.slm", `DDR_X_BRAM_RAMLOOP(187) );
  $readmemh("slm_files/ddr_x_mem_cut28_5.slm", `DDR_X_BRAM_RAMLOOP(188) );
  $readmemh("slm_files/ddr_x_mem_cut29_5.slm", `DDR_X_BRAM_RAMLOOP(189) );
  $readmemh("slm_files/ddr_x_mem_cut30_5.slm", `DDR_X_BRAM_RAMLOOP(190) );
  $readmemh("slm_files/ddr_x_mem_cut31_5.slm", `DDR_X_BRAM_RAMLOOP(191) );
  $readmemh("slm_files/ddr_x_mem_cut0_6.slm", `DDR_X_BRAM_RAMLOOP(192) );
  $readmemh("slm_files/ddr_x_mem_cut1_6.slm", `DDR_X_BRAM_RAMLOOP(193) );
  $readmemh("slm_files/ddr_x_mem_cut2_6.slm", `DDR_X_BRAM_RAMLOOP(194) );
  $readmemh("slm_files/ddr_x_mem_cut3_6.slm", `DDR_X_BRAM_RAMLOOP(195) );
  $readmemh("slm_files/ddr_x_mem_cut4_6.slm", `DDR_X_BRAM_RAMLOOP(196) );
  $readmemh("slm_files/ddr_x_mem_cut5_6.slm", `DDR_X_BRAM_RAMLOOP(197) );
  $readmemh("slm_files/ddr_x_mem_cut6_6.slm", `DDR_X_BRAM_RAMLOOP(198) );
  $readmemh("slm_files/ddr_x_mem_cut7_6.slm", `DDR_X_BRAM_RAMLOOP(199) );
  $readmemh("slm_files/ddr_x_mem_cut8_6.slm", `DDR_X_BRAM_RAMLOOP(200) );
  $readmemh("slm_files/ddr_x_mem_cut9_6.slm", `DDR_X_BRAM_RAMLOOP(201) );
  $readmemh("slm_files/ddr_x_mem_cut10_6.slm", `DDR_X_BRAM_RAMLOOP(202) );
  $readmemh("slm_files/ddr_x_mem_cut11_6.slm", `DDR_X_BRAM_RAMLOOP(203) );
  $readmemh("slm_files/ddr_x_mem_cut12_6.slm", `DDR_X_BRAM_RAMLOOP(204) );
  $readmemh("slm_files/ddr_x_mem_cut13_6.slm", `DDR_X_BRAM_RAMLOOP(205) );
  $readmemh("slm_files/ddr_x_mem_cut14_6.slm", `DDR_X_BRAM_RAMLOOP(206) );
  $readmemh("slm_files/ddr_x_mem_cut15_6.slm", `DDR_X_BRAM_RAMLOOP(207) );
  $readmemh("slm_files/ddr_x_mem_cut16_6.slm", `DDR_X_BRAM_RAMLOOP(208) );
  $readmemh("slm_files/ddr_x_mem_cut17_6.slm", `DDR_X_BRAM_RAMLOOP(209) );
  $readmemh("slm_files/ddr_x_mem_cut18_6.slm", `DDR_X_BRAM_RAMLOOP(210) );
  $readmemh("slm_files/ddr_x_mem_cut19_6.slm", `DDR_X_BRAM_RAMLOOP(211) );
  $readmemh("slm_files/ddr_x_mem_cut20_6.slm", `DDR_X_BRAM_RAMLOOP(212) );
  $readmemh("slm_files/ddr_x_mem_cut21_6.slm", `DDR_X_BRAM_RAMLOOP(213) );
  $readmemh("slm_files/ddr_x_mem_cut22_6.slm", `DDR_X_BRAM_RAMLOOP(214) );
  $readmemh("slm_files/ddr_x_mem_cut23_6.slm", `DDR_X_BRAM_RAMLOOP(215) );
  $readmemh("slm_files/ddr_x_mem_cut24_6.slm", `DDR_X_BRAM_RAMLOOP(216) );
  $readmemh("slm_files/ddr_x_mem_cut25_6.slm", `DDR_X_BRAM_RAMLOOP(217) );
  $readmemh("slm_files/ddr_x_mem_cut26_6.slm", `DDR_X_BRAM_RAMLOOP(218) );
  $readmemh("slm_files/ddr_x_mem_cut27_6.slm", `DDR_X_BRAM_RAMLOOP(219) );
  $readmemh("slm_files/ddr_x_mem_cut28_6.slm", `DDR_X_BRAM_RAMLOOP(220) );
  $readmemh("slm_files/ddr_x_mem_cut29_6.slm", `DDR_X_BRAM_RAMLOOP(221) );
  $readmemh("slm_files/ddr_x_mem_cut30_6.slm", `DDR_X_BRAM_RAMLOOP(222) );
  $readmemh("slm_files/ddr_x_mem_cut31_6.slm", `DDR_X_BRAM_RAMLOOP(223) );
  $readmemh("slm_files/ddr_x_mem_cut0_7.slm", `DDR_X_BRAM_RAMLOOP(224) );
  $readmemh("slm_files/ddr_x_mem_cut1_7.slm", `DDR_X_BRAM_RAMLOOP(225) );
  $readmemh("slm_files/ddr_x_mem_cut2_7.slm", `DDR_X_BRAM_RAMLOOP(226) );
  $readmemh("slm_files/ddr_x_mem_cut3_7.slm", `DDR_X_BRAM_RAMLOOP(227) );
  $readmemh("slm_files/ddr_x_mem_cut4_7.slm", `DDR_X_BRAM_RAMLOOP(228) );
  $readmemh("slm_files/ddr_x_mem_cut5_7.slm", `DDR_X_BRAM_RAMLOOP(229) );
  $readmemh("slm_files/ddr_x_mem_cut6_7.slm", `DDR_X_BRAM_RAMLOOP(230) );
  $readmemh("slm_files/ddr_x_mem_cut7_7.slm", `DDR_X_BRAM_RAMLOOP(231) );
  $readmemh("slm_files/ddr_x_mem_cut8_7.slm", `DDR_X_BRAM_RAMLOOP(232) );
  $readmemh("slm_files/ddr_x_mem_cut9_7.slm", `DDR_X_BRAM_RAMLOOP(233) );
  $readmemh("slm_files/ddr_x_mem_cut10_7.slm", `DDR_X_BRAM_RAMLOOP(234) );
  $readmemh("slm_files/ddr_x_mem_cut11_7.slm", `DDR_X_BRAM_RAMLOOP(235) );
  $readmemh("slm_files/ddr_x_mem_cut12_7.slm", `DDR_X_BRAM_RAMLOOP(236) );
  $readmemh("slm_files/ddr_x_mem_cut13_7.slm", `DDR_X_BRAM_RAMLOOP(237) );
  $readmemh("slm_files/ddr_x_mem_cut14_7.slm", `DDR_X_BRAM_RAMLOOP(238) );
  $readmemh("slm_files/ddr_x_mem_cut15_7.slm", `DDR_X_BRAM_RAMLOOP(239) );
  $readmemh("slm_files/ddr_x_mem_cut16_7.slm", `DDR_X_BRAM_RAMLOOP(240) );
  $readmemh("slm_files/ddr_x_mem_cut17_7.slm", `DDR_X_BRAM_RAMLOOP(241) );
  $readmemh("slm_files/ddr_x_mem_cut18_7.slm", `DDR_X_BRAM_RAMLOOP(242) );
  $readmemh("slm_files/ddr_x_mem_cut19_7.slm", `DDR_X_BRAM_RAMLOOP(243) );
  $readmemh("slm_files/ddr_x_mem_cut20_7.slm", `DDR_X_BRAM_RAMLOOP(244) );
  $readmemh("slm_files/ddr_x_mem_cut21_7.slm", `DDR_X_BRAM_RAMLOOP(245) );
  $readmemh("slm_files/ddr_x_mem_cut22_7.slm", `DDR_X_BRAM_RAMLOOP(246) );
  $readmemh("slm_files/ddr_x_mem_cut23_7.slm", `DDR_X_BRAM_RAMLOOP(247) );
  $readmemh("slm_files/ddr_x_mem_cut24_7.slm", `DDR_X_BRAM_RAMLOOP(248) );
  $readmemh("slm_files/ddr_x_mem_cut25_7.slm", `DDR_X_BRAM_RAMLOOP(249) );
  $readmemh("slm_files/ddr_x_mem_cut26_7.slm", `DDR_X_BRAM_RAMLOOP(250) );
  $readmemh("slm_files/ddr_x_mem_cut27_7.slm", `DDR_X_BRAM_RAMLOOP(251) );
  $readmemh("slm_files/ddr_x_mem_cut28_7.slm", `DDR_X_BRAM_RAMLOOP(252) );
  $readmemh("slm_files/ddr_x_mem_cut29_7.slm", `DDR_X_BRAM_RAMLOOP(253) );
  $readmemh("slm_files/ddr_x_mem_cut30_7.slm", `DDR_X_BRAM_RAMLOOP(254) );
  $readmemh("slm_files/ddr_x_mem_cut31_7.slm", `DDR_X_BRAM_RAMLOOP(255) );
endtask
